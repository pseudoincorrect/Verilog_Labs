library verilog;
use verilog.vl_types.all;
entity mesh_testbench is
end mesh_testbench;
