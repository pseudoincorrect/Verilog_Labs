library verilog;
use verilog.vl_types.all;
entity node_testbench is
end node_testbench;
