-- megafunction wizard: %ALTFP_MULT%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: ALTFP_MULT 

-- ============================================================
-- File Name: mult.vhd
-- Megafunction Name(s):
-- 			ALTFP_MULT
--
-- Simulation Library Files(s):
-- 			lpm
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 13.0.1 Build 232 06/12/2013 SP 1 SJ Web Edition
-- ************************************************************


--Copyright (C) 1991-2013 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


--altfp_mult CBX_AUTO_BLACKBOX="ALL" DEDICATED_MULTIPLIER_CIRCUITRY="YES" DENORMAL_SUPPORT="NO" DEVICE_FAMILY="Cyclone IV GX" EXCEPTION_HANDLING="NO" PIPELINE=5 REDUCED_FUNCTIONALITY="NO" ROUNDING="TO_NEAREST" WIDTH_EXP=11 WIDTH_MAN=52 clock dataa datab overflow result
--VERSION_BEGIN 13.0 cbx_alt_ded_mult_y 2013:06:12:18:03:43:SJ cbx_altbarrel_shift 2013:06:12:18:03:43:SJ cbx_altera_mult_add 2013:06:12:18:03:43:SJ cbx_altera_mult_add_rtl 2013:06:12:18:03:43:SJ cbx_altfp_mult 2013:06:12:18:03:43:SJ cbx_altmult_add 2013:06:12:18:03:43:SJ cbx_cycloneii 2013:06:12:18:03:43:SJ cbx_lpm_add_sub 2013:06:12:18:03:43:SJ cbx_lpm_compare 2013:06:12:18:03:43:SJ cbx_lpm_mult 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ cbx_padd 2013:06:12:18:03:43:SJ cbx_parallel_add 2013:06:12:18:03:43:SJ cbx_stratix 2013:06:12:18:03:43:SJ cbx_stratixii 2013:06:12:18:03:43:SJ cbx_util_mgl 2013:06:12:18:03:43:SJ  VERSION_END

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = lpm_add_sub 4 lpm_mult 1 reg 236 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  mult_altfp_mult_nto IS 
	 PORT 
	 ( 
		 clock	:	IN  STD_LOGIC;
		 dataa	:	IN  STD_LOGIC_VECTOR (63 DOWNTO 0);
		 datab	:	IN  STD_LOGIC_VECTOR (63 DOWNTO 0);
		 overflow	:	OUT  STD_LOGIC;
		 result	:	OUT  STD_LOGIC_VECTOR (63 DOWNTO 0)
	 ); 
 END mult_altfp_mult_nto;

 ARCHITECTURE RTL OF mult_altfp_mult_nto IS

	 SIGNAL	 dataa_exp_all_one_ff_p1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_dataa_exp_all_one_ff_p1_w_lg_q512w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dataa_exp_all_one_ff_p1_w_lg_q507w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 dataa_exp_not_zero_ff_p1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 dataa_man_not_zero_ff_p1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_dataa_man_not_zero_ff_p1_w_lg_w_lg_q506w511w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dataa_man_not_zero_ff_p1_w_lg_q506w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 dataa_man_not_zero_ff_p2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 datab_exp_all_one_ff_p1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_datab_exp_all_one_ff_p1_w_lg_q510w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_datab_exp_all_one_ff_p1_w_lg_q505w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 datab_exp_not_zero_ff_p1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 datab_man_not_zero_ff_p1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_datab_man_not_zero_ff_p1_w_lg_w_lg_q504w509w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_datab_man_not_zero_ff_p1_w_lg_q504w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 datab_man_not_zero_ff_p2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 delay_exp2_bias	:	STD_LOGIC_VECTOR(12 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 delay_exp_bias	:	STD_LOGIC_VECTOR(12 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 delay_man_product_msb	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_delay_man_product_msb_w_lg_q696w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_delay_man_product_msb_w_lg_q698w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 delay_man_product_msb_p0	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_add_p1	:	STD_LOGIC_VECTOR(11 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_result_ff	:	STD_LOGIC_VECTOR(10 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_dffe_0	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_dffe_1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_ff1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_input_is_infinity_ff1_w_lg_q780w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_input_is_infinity_ff1_w_lg_q786w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 input_is_nan_dffe_0	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_dffe_1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_ff1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_input_is_nan_ff1_w_lg_q782w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 input_not_zero_dffe_0	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_not_zero_dffe_1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_not_zero_ff1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_input_not_zero_ff1_w_lg_q779w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 lsb_dffe	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 man_result_ff	:	STD_LOGIC_VECTOR(51 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 man_round_p	:	STD_LOGIC_VECTOR(52 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 man_round_p2	:	STD_LOGIC_VECTOR(53 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_man_round_p2_w_lg_w_q_range702w703w	:	STD_LOGIC_VECTOR (52 DOWNTO 0);
	 SIGNAL  wire_man_round_p2_w_lg_w_q_range699w700w	:	STD_LOGIC_VECTOR (52 DOWNTO 0);
	 SIGNAL  wire_man_round_p2_w_lg_w_q_range694w701w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_round_p2_w_q_range702w	:	STD_LOGIC_VECTOR (52 DOWNTO 0);
	 SIGNAL  wire_man_round_p2_w_q_range699w	:	STD_LOGIC_VECTOR (52 DOWNTO 0);
	 SIGNAL  wire_man_round_p2_w_q_range694w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 overflow_ff	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 round_dffe	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_node_ff0	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_node_ff1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_node_ff2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_node_ff3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_node_ff4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sticky_dffe	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_gnd	:	STD_LOGIC;
	 SIGNAL  wire_exp_add_adder_dataa	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  wire_exp_add_adder_datab	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  wire_exp_add_adder_result	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  wire_exp_adj_adder_w_lg_w_lg_w_result_range772w773w774w	:	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  wire_exp_adj_adder_w_lg_w_result_range772w773w	:	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  wire_exp_adj_adder_w_lg_w_result_range739w770w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_adj_adder_result	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_exp_adj_adder_w_result_range772w	:	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  wire_exp_adj_adder_w_result_range735w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_adj_adder_w_result_range738w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_adj_adder_w_result_range739w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_adj_adder_w_result_range708w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_adj_adder_w_result_range711w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_adj_adder_w_result_range714w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_adj_adder_w_result_range717w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_adj_adder_w_result_range720w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_adj_adder_w_result_range723w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_adj_adder_w_result_range726w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_adj_adder_w_result_range729w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_adj_adder_w_result_range732w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_bias_subtr_dataa	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_exp_bias_subtr_datab	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_exp_bias_subtr_result	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_man_round_adder_dataa	:	STD_LOGIC_VECTOR (53 DOWNTO 0);
	 SIGNAL  wire_man_round_adder_datab	:	STD_LOGIC_VECTOR (53 DOWNTO 0);
	 SIGNAL  wire_man_round_adder_result	:	STD_LOGIC_VECTOR (53 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_lg_w_result_range518w519w	:	STD_LOGIC_VECTOR (53 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_lg_w_result_range514w676w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_lg_w_result_range515w516w	:	STD_LOGIC_VECTOR (53 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_lg_w_result_range514w517w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_dataa	:	STD_LOGIC_VECTOR (52 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_datab	:	STD_LOGIC_VECTOR (52 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_result	:	STD_LOGIC_VECTOR (105 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range518w	:	STD_LOGIC_VECTOR (53 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range514w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range515w	:	STD_LOGIC_VECTOR (53 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range551w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range554w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range557w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range560w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range563w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range566w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range569w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range572w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range575w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range578w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range524w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range581w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range584w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range587w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range590w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range593w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range596w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range599w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range602w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range605w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range608w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range527w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range611w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range614w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range617w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range620w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range623w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range626w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range629w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range632w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range635w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range638w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range530w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range641w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range644w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range647w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range650w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range653w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range656w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range659w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range662w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range665w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range668w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range533w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range671w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range674w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range536w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range539w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range542w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range545w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range548w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w799w800w801w	:	STD_LOGIC_VECTOR (50 DOWNTO 0);
	 SIGNAL  wire_w_lg_w799w800w	:	STD_LOGIC_VECTOR (50 DOWNTO 0);
	 SIGNAL  wire_w_lg_w790w791w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w799w	:	STD_LOGIC_VECTOR (50 DOWNTO 0);
	 SIGNAL  wire_w790w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_man_result_round_range796w797w798w	:	STD_LOGIC_VECTOR (50 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_man_result_round_range787w788w789w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_inf_num777w	:	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range93w100w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range103w110w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range113w120w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range123w130w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range133w140w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range143w150w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range153w160w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range163w170w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range173w180w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range183w190w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range96w102w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range106w112w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range116w122w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range126w132w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range136w142w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range146w152w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range156w162w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range166w172w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range176w182w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range186w192w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_result_round_range796w797w	:	STD_LOGIC_VECTOR (50 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_result_round_range787w788w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_result_exp_all_one_range706w710w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_result_exp_all_one_range709w713w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_result_exp_all_one_range712w716w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_result_exp_all_one_range715w719w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_result_exp_all_one_range718w722w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_result_exp_all_one_range721w725w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_result_exp_all_one_range724w728w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_result_exp_all_one_range727w731w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_result_exp_all_one_range730w734w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_result_exp_all_one_range733w737w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_exp_is_inf785w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_exp_is_zero771w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_result_exp_not_zero_range767w769w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w790w791w792w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_inf_num777w778w	:	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w790w791w792w793w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_exp_is_inf775w776w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_exp_is_inf775w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range253w255w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range259w261w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range265w267w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range271w273w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range277w279w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range283w285w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range289w291w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range295w297w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range301w303w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range307w309w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range199w201w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range313w315w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range319w321w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range325w327w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range331w333w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range337w339w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range343w345w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range353w355w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range359w361w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range365w367w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range205w207w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range371w373w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range377w379w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range383w385w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range389w391w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range395w397w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range401w403w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range407w409w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range413w415w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range419w421w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range425w427w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range211w213w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range431w433w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range437w439w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range443w445w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range449w451w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range455w457w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range461w463w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range467w469w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range473w475w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range479w481w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range485w487w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range217w219w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range491w493w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range497w499w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range93w95w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range103w105w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range113w115w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range123w125w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range133w135w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range143w145w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range153w155w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range223w225w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range163w165w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range173w175w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range183w185w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range229w231w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range235w237w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range241w243w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range247w249w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range256w258w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range262w264w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range268w270w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range274w276w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range280w282w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range286w288w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range292w294w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range298w300w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range304w306w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range310w312w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range202w204w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range316w318w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range322w324w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range328w330w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range334w336w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range340w342w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range346w348w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range356w358w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range362w364w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range368w370w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range208w210w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range374w376w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range380w382w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range386w388w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range392w394w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range398w400w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range404w406w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range410w412w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range416w418w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range422w424w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range428w430w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range214w216w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range434w436w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range440w442w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range446w448w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range452w454w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range458w460w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range464w466w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range470w472w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range476w478w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range482w484w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range488w490w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range220w222w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range494w496w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range500w502w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range96w98w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range106w108w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range116w118w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range126w128w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range136w138w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range146w148w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range156w158w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range226w228w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range166w168w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range176w178w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range186w188w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range232w234w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range238w240w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range244w246w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range250w252w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_result_exp_not_zero_range745w748w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_result_exp_not_zero_range765w768w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_result_exp_not_zero_range747w750w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_result_exp_not_zero_range749w752w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_result_exp_not_zero_range751w754w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_result_exp_not_zero_range753w756w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_result_exp_not_zero_range755w758w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_result_exp_not_zero_range757w760w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_result_exp_not_zero_range759w762w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_result_exp_not_zero_range761w764w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_result_exp_not_zero_range763w766w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_range522w526w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_range552w556w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_range555w559w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_range558w562w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_range561w565w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_range564w568w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_range567w571w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_range570w574w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_range573w577w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_range576w580w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_range579w583w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_range525w529w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_range582w586w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_range585w589w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_range588w592w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_range591w595w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_range594w598w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_range597w601w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_range600w604w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_range603w607w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_range606w610w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_range609w613w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_range528w532w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_range612w616w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_range615w619w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_range618w622w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_range621w625w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_range624w628w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_range627w631w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_range630w634w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_range633w637w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_range636w640w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_range639w643w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_range531w535w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_range642w646w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_range645w649w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_range648w652w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_range651w655w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_range654w658w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_range657w661w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_range660w664w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_range663w667w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_range666w670w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_range669w673w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_range534w538w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_range672w677w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_range537w541w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_range540w544w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_range543w547w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_range546w550w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_range549w553w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  aclr	:	STD_LOGIC;
	 SIGNAL  bias :	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  clk_en	:	STD_LOGIC;
	 SIGNAL  dataa_exp_all_one :	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  dataa_exp_not_zero :	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  dataa_man_not_zero :	STD_LOGIC_VECTOR (51 DOWNTO 0);
	 SIGNAL  datab_exp_all_one :	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  datab_exp_not_zero :	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  datab_man_not_zero :	STD_LOGIC_VECTOR (51 DOWNTO 0);
	 SIGNAL  exp_is_inf :	STD_LOGIC;
	 SIGNAL  exp_is_zero :	STD_LOGIC;
	 SIGNAL  expmod :	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  inf_num :	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  lsb_bit :	STD_LOGIC;
	 SIGNAL  man_result_round :	STD_LOGIC_VECTOR (52 DOWNTO 0);
	 SIGNAL  man_shift_full :	STD_LOGIC_VECTOR (53 DOWNTO 0);
	 SIGNAL  result_exp_all_one :	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  result_exp_not_zero :	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  round_bit :	STD_LOGIC;
	 SIGNAL  round_carry :	STD_LOGIC;
	 SIGNAL  sticky_bit :	STD_LOGIC_VECTOR (51 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range253w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range259w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range265w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range271w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range277w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range283w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range289w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range295w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range301w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range307w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range199w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range313w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range319w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range325w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range331w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range337w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range343w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range353w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range359w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range365w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range205w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range371w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range377w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range383w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range389w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range395w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range401w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range407w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range413w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range419w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range425w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range211w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range431w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range437w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range443w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range449w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range455w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range461w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range467w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range473w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range479w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range485w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range217w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range491w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range497w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range93w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range103w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range113w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range123w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range133w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range143w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range153w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range223w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range163w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range173w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range183w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range229w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range235w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range241w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range247w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_exp_all_one_range89w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_exp_all_one_range99w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_exp_all_one_range109w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_exp_all_one_range119w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_exp_all_one_range129w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_exp_all_one_range139w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_exp_all_one_range149w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_exp_all_one_range159w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_exp_all_one_range169w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_exp_all_one_range179w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_exp_not_zero_range84w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_exp_not_zero_range94w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_exp_not_zero_range104w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_exp_not_zero_range114w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_exp_not_zero_range124w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_exp_not_zero_range134w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_exp_not_zero_range144w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_exp_not_zero_range154w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_exp_not_zero_range164w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_exp_not_zero_range174w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_man_not_zero_range194w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_man_not_zero_range254w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_man_not_zero_range260w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_man_not_zero_range266w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_man_not_zero_range272w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_man_not_zero_range278w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_man_not_zero_range284w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_man_not_zero_range290w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_man_not_zero_range296w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_man_not_zero_range302w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_man_not_zero_range308w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_man_not_zero_range200w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_man_not_zero_range314w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_man_not_zero_range320w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_man_not_zero_range326w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_man_not_zero_range332w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_man_not_zero_range338w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_man_not_zero_range350w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_man_not_zero_range354w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_man_not_zero_range360w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_man_not_zero_range366w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_man_not_zero_range206w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_man_not_zero_range372w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_man_not_zero_range378w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_man_not_zero_range384w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_man_not_zero_range390w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_man_not_zero_range396w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_man_not_zero_range402w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_man_not_zero_range408w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_man_not_zero_range414w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_man_not_zero_range420w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_man_not_zero_range426w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_man_not_zero_range212w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_man_not_zero_range432w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_man_not_zero_range438w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_man_not_zero_range444w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_man_not_zero_range450w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_man_not_zero_range456w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_man_not_zero_range462w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_man_not_zero_range468w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_man_not_zero_range474w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_man_not_zero_range480w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_man_not_zero_range486w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_man_not_zero_range218w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_man_not_zero_range492w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_man_not_zero_range224w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_man_not_zero_range230w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_man_not_zero_range236w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_man_not_zero_range242w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_man_not_zero_range248w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range256w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range262w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range268w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range274w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range280w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range286w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range292w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range298w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range304w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range310w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range202w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range316w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range322w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range328w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range334w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range340w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range346w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range356w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range362w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range368w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range208w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range374w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range380w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range386w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range392w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range398w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range404w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range410w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range416w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range422w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range428w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range214w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range434w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range440w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range446w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range452w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range458w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range464w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range470w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range476w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range482w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range488w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range220w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range494w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range500w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range96w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range106w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range116w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range126w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range136w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range146w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range156w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range226w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range166w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range176w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range186w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range232w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range238w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range244w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range250w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_exp_all_one_range91w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_exp_all_one_range101w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_exp_all_one_range111w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_exp_all_one_range121w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_exp_all_one_range131w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_exp_all_one_range141w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_exp_all_one_range151w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_exp_all_one_range161w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_exp_all_one_range171w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_exp_all_one_range181w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_exp_not_zero_range87w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_exp_not_zero_range97w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_exp_not_zero_range107w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_exp_not_zero_range117w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_exp_not_zero_range127w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_exp_not_zero_range137w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_exp_not_zero_range147w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_exp_not_zero_range157w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_exp_not_zero_range167w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_exp_not_zero_range177w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_man_not_zero_range197w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_man_not_zero_range257w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_man_not_zero_range263w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_man_not_zero_range269w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_man_not_zero_range275w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_man_not_zero_range281w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_man_not_zero_range287w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_man_not_zero_range293w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_man_not_zero_range299w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_man_not_zero_range305w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_man_not_zero_range311w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_man_not_zero_range203w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_man_not_zero_range317w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_man_not_zero_range323w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_man_not_zero_range329w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_man_not_zero_range335w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_man_not_zero_range341w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_man_not_zero_range352w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_man_not_zero_range357w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_man_not_zero_range363w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_man_not_zero_range369w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_man_not_zero_range209w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_man_not_zero_range375w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_man_not_zero_range381w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_man_not_zero_range387w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_man_not_zero_range393w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_man_not_zero_range399w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_man_not_zero_range405w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_man_not_zero_range411w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_man_not_zero_range417w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_man_not_zero_range423w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_man_not_zero_range429w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_man_not_zero_range215w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_man_not_zero_range435w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_man_not_zero_range441w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_man_not_zero_range447w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_man_not_zero_range453w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_man_not_zero_range459w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_man_not_zero_range465w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_man_not_zero_range471w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_man_not_zero_range477w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_man_not_zero_range483w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_man_not_zero_range489w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_man_not_zero_range221w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_man_not_zero_range495w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_man_not_zero_range227w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_man_not_zero_range233w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_man_not_zero_range239w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_man_not_zero_range245w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_man_not_zero_range251w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_result_round_range796w	:	STD_LOGIC_VECTOR (50 DOWNTO 0);
	 SIGNAL  wire_w_man_result_round_range787w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_shift_full_range682w	:	STD_LOGIC_VECTOR (52 DOWNTO 0);
	 SIGNAL  wire_w_result_exp_all_one_range706w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_result_exp_all_one_range709w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_result_exp_all_one_range712w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_result_exp_all_one_range715w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_result_exp_all_one_range718w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_result_exp_all_one_range721w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_result_exp_all_one_range724w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_result_exp_all_one_range727w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_result_exp_all_one_range730w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_result_exp_all_one_range733w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_result_exp_not_zero_range745w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_result_exp_not_zero_range765w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_result_exp_not_zero_range767w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_result_exp_not_zero_range747w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_result_exp_not_zero_range749w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_result_exp_not_zero_range751w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_result_exp_not_zero_range753w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_result_exp_not_zero_range755w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_result_exp_not_zero_range757w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_result_exp_not_zero_range759w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_result_exp_not_zero_range761w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_result_exp_not_zero_range763w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_range522w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_range552w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_range555w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_range558w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_range561w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_range564w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_range567w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_range570w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_range573w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_range576w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_range579w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_range525w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_range582w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_range585w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_range588w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_range591w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_range594w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_range597w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_range600w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_range603w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_range606w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_range609w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_range528w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_range612w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_range615w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_range618w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_range621w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_range624w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_range627w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_range630w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_range633w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_range636w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_range639w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_range531w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_range642w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_range645w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_range648w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_range651w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_range654w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_range657w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_range660w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_range663w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_range666w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_range669w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_range534w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_range672w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_range537w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_range540w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_range543w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_range546w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_range549w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_mult
	 GENERIC 
	 (
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "UNSIGNED";
		LPM_WIDTHA	:	NATURAL;
		LPM_WIDTHB	:	NATURAL;
		LPM_WIDTHP	:	NATURAL;
		LPM_WIDTHS	:	NATURAL := 1;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_mult"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTHA-1 DOWNTO 0);
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTHB-1 DOWNTO 0);
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTHP-1 DOWNTO 0);
		sum	:	IN STD_LOGIC_VECTOR(LPM_WIDTHS-1 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
 BEGIN

	wire_gnd <= '0';
	loop0 : FOR i IN 0 TO 50 GENERATE 
		wire_w_lg_w_lg_w799w800w801w(i) <= wire_w_lg_w799w800w(i) AND wire_input_is_nan_ff1_w_lg_q782w(0);
	END GENERATE loop0;
	loop1 : FOR i IN 0 TO 50 GENERATE 
		wire_w_lg_w799w800w(i) <= wire_w799w(i) AND wire_w_lg_exp_is_zero771w(0);
	END GENERATE loop1;
	wire_w_lg_w790w791w(0) <= wire_w790w(0) AND wire_w_lg_exp_is_zero771w(0);
	loop2 : FOR i IN 0 TO 50 GENERATE 
		wire_w799w(i) <= wire_w_lg_w_lg_w_man_result_round_range796w797w798w(i) AND wire_w_lg_exp_is_inf785w(0);
	END GENERATE loop2;
	wire_w790w(0) <= wire_w_lg_w_lg_w_man_result_round_range787w788w789w(0) AND wire_w_lg_exp_is_inf785w(0);
	loop3 : FOR i IN 0 TO 50 GENERATE 
		wire_w_lg_w_lg_w_man_result_round_range796w797w798w(i) <= wire_w_lg_w_man_result_round_range796w797w(i) AND wire_input_is_infinity_ff1_w_lg_q786w(0);
	END GENERATE loop3;
	wire_w_lg_w_lg_w_man_result_round_range787w788w789w(0) <= wire_w_lg_w_man_result_round_range787w788w(0) AND wire_input_is_infinity_ff1_w_lg_q786w(0);
	loop4 : FOR i IN 0 TO 10 GENERATE 
		wire_w_lg_inf_num777w(i) <= inf_num(i) AND wire_w_lg_w_lg_exp_is_inf775w776w(0);
	END GENERATE loop4;
	wire_w_lg_w_dataa_range93w100w(0) <= wire_w_dataa_range93w(0) AND wire_w_dataa_exp_all_one_range89w(0);
	wire_w_lg_w_dataa_range103w110w(0) <= wire_w_dataa_range103w(0) AND wire_w_dataa_exp_all_one_range99w(0);
	wire_w_lg_w_dataa_range113w120w(0) <= wire_w_dataa_range113w(0) AND wire_w_dataa_exp_all_one_range109w(0);
	wire_w_lg_w_dataa_range123w130w(0) <= wire_w_dataa_range123w(0) AND wire_w_dataa_exp_all_one_range119w(0);
	wire_w_lg_w_dataa_range133w140w(0) <= wire_w_dataa_range133w(0) AND wire_w_dataa_exp_all_one_range129w(0);
	wire_w_lg_w_dataa_range143w150w(0) <= wire_w_dataa_range143w(0) AND wire_w_dataa_exp_all_one_range139w(0);
	wire_w_lg_w_dataa_range153w160w(0) <= wire_w_dataa_range153w(0) AND wire_w_dataa_exp_all_one_range149w(0);
	wire_w_lg_w_dataa_range163w170w(0) <= wire_w_dataa_range163w(0) AND wire_w_dataa_exp_all_one_range159w(0);
	wire_w_lg_w_dataa_range173w180w(0) <= wire_w_dataa_range173w(0) AND wire_w_dataa_exp_all_one_range169w(0);
	wire_w_lg_w_dataa_range183w190w(0) <= wire_w_dataa_range183w(0) AND wire_w_dataa_exp_all_one_range179w(0);
	wire_w_lg_w_datab_range96w102w(0) <= wire_w_datab_range96w(0) AND wire_w_datab_exp_all_one_range91w(0);
	wire_w_lg_w_datab_range106w112w(0) <= wire_w_datab_range106w(0) AND wire_w_datab_exp_all_one_range101w(0);
	wire_w_lg_w_datab_range116w122w(0) <= wire_w_datab_range116w(0) AND wire_w_datab_exp_all_one_range111w(0);
	wire_w_lg_w_datab_range126w132w(0) <= wire_w_datab_range126w(0) AND wire_w_datab_exp_all_one_range121w(0);
	wire_w_lg_w_datab_range136w142w(0) <= wire_w_datab_range136w(0) AND wire_w_datab_exp_all_one_range131w(0);
	wire_w_lg_w_datab_range146w152w(0) <= wire_w_datab_range146w(0) AND wire_w_datab_exp_all_one_range141w(0);
	wire_w_lg_w_datab_range156w162w(0) <= wire_w_datab_range156w(0) AND wire_w_datab_exp_all_one_range151w(0);
	wire_w_lg_w_datab_range166w172w(0) <= wire_w_datab_range166w(0) AND wire_w_datab_exp_all_one_range161w(0);
	wire_w_lg_w_datab_range176w182w(0) <= wire_w_datab_range176w(0) AND wire_w_datab_exp_all_one_range171w(0);
	wire_w_lg_w_datab_range186w192w(0) <= wire_w_datab_range186w(0) AND wire_w_datab_exp_all_one_range181w(0);
	loop5 : FOR i IN 0 TO 50 GENERATE 
		wire_w_lg_w_man_result_round_range796w797w(i) <= wire_w_man_result_round_range796w(i) AND input_not_zero_ff1;
	END GENERATE loop5;
	wire_w_lg_w_man_result_round_range787w788w(0) <= wire_w_man_result_round_range787w(0) AND input_not_zero_ff1;
	wire_w_lg_w_result_exp_all_one_range706w710w(0) <= wire_w_result_exp_all_one_range706w(0) AND wire_exp_adj_adder_w_result_range708w(0);
	wire_w_lg_w_result_exp_all_one_range709w713w(0) <= wire_w_result_exp_all_one_range709w(0) AND wire_exp_adj_adder_w_result_range711w(0);
	wire_w_lg_w_result_exp_all_one_range712w716w(0) <= wire_w_result_exp_all_one_range712w(0) AND wire_exp_adj_adder_w_result_range714w(0);
	wire_w_lg_w_result_exp_all_one_range715w719w(0) <= wire_w_result_exp_all_one_range715w(0) AND wire_exp_adj_adder_w_result_range717w(0);
	wire_w_lg_w_result_exp_all_one_range718w722w(0) <= wire_w_result_exp_all_one_range718w(0) AND wire_exp_adj_adder_w_result_range720w(0);
	wire_w_lg_w_result_exp_all_one_range721w725w(0) <= wire_w_result_exp_all_one_range721w(0) AND wire_exp_adj_adder_w_result_range723w(0);
	wire_w_lg_w_result_exp_all_one_range724w728w(0) <= wire_w_result_exp_all_one_range724w(0) AND wire_exp_adj_adder_w_result_range726w(0);
	wire_w_lg_w_result_exp_all_one_range727w731w(0) <= wire_w_result_exp_all_one_range727w(0) AND wire_exp_adj_adder_w_result_range729w(0);
	wire_w_lg_w_result_exp_all_one_range730w734w(0) <= wire_w_result_exp_all_one_range730w(0) AND wire_exp_adj_adder_w_result_range732w(0);
	wire_w_lg_w_result_exp_all_one_range733w737w(0) <= wire_w_result_exp_all_one_range733w(0) AND wire_exp_adj_adder_w_result_range735w(0);
	wire_w_lg_exp_is_inf785w(0) <= NOT exp_is_inf;
	wire_w_lg_exp_is_zero771w(0) <= NOT exp_is_zero;
	wire_w_lg_w_result_exp_not_zero_range767w769w(0) <= NOT wire_w_result_exp_not_zero_range767w(0);
	wire_w_lg_w_lg_w790w791w792w(0) <= wire_w_lg_w790w791w(0) OR wire_input_is_infinity_ff1_w_lg_q780w(0);
	loop6 : FOR i IN 0 TO 10 GENERATE 
		wire_w_lg_w_lg_inf_num777w778w(i) <= wire_w_lg_inf_num777w(i) OR wire_exp_adj_adder_w_lg_w_lg_w_result_range772w773w774w(i);
	END GENERATE loop6;
	wire_w_lg_w_lg_w_lg_w790w791w792w793w(0) <= wire_w_lg_w_lg_w790w791w792w(0) OR input_is_nan_ff1;
	wire_w_lg_w_lg_exp_is_inf775w776w(0) <= wire_w_lg_exp_is_inf775w(0) OR input_is_nan_ff1;
	wire_w_lg_exp_is_inf775w(0) <= exp_is_inf OR input_is_infinity_ff1;
	wire_w_lg_w_dataa_range253w255w(0) <= wire_w_dataa_range253w(0) OR wire_w_dataa_man_not_zero_range248w(0);
	wire_w_lg_w_dataa_range259w261w(0) <= wire_w_dataa_range259w(0) OR wire_w_dataa_man_not_zero_range254w(0);
	wire_w_lg_w_dataa_range265w267w(0) <= wire_w_dataa_range265w(0) OR wire_w_dataa_man_not_zero_range260w(0);
	wire_w_lg_w_dataa_range271w273w(0) <= wire_w_dataa_range271w(0) OR wire_w_dataa_man_not_zero_range266w(0);
	wire_w_lg_w_dataa_range277w279w(0) <= wire_w_dataa_range277w(0) OR wire_w_dataa_man_not_zero_range272w(0);
	wire_w_lg_w_dataa_range283w285w(0) <= wire_w_dataa_range283w(0) OR wire_w_dataa_man_not_zero_range278w(0);
	wire_w_lg_w_dataa_range289w291w(0) <= wire_w_dataa_range289w(0) OR wire_w_dataa_man_not_zero_range284w(0);
	wire_w_lg_w_dataa_range295w297w(0) <= wire_w_dataa_range295w(0) OR wire_w_dataa_man_not_zero_range290w(0);
	wire_w_lg_w_dataa_range301w303w(0) <= wire_w_dataa_range301w(0) OR wire_w_dataa_man_not_zero_range296w(0);
	wire_w_lg_w_dataa_range307w309w(0) <= wire_w_dataa_range307w(0) OR wire_w_dataa_man_not_zero_range302w(0);
	wire_w_lg_w_dataa_range199w201w(0) <= wire_w_dataa_range199w(0) OR wire_w_dataa_man_not_zero_range194w(0);
	wire_w_lg_w_dataa_range313w315w(0) <= wire_w_dataa_range313w(0) OR wire_w_dataa_man_not_zero_range308w(0);
	wire_w_lg_w_dataa_range319w321w(0) <= wire_w_dataa_range319w(0) OR wire_w_dataa_man_not_zero_range314w(0);
	wire_w_lg_w_dataa_range325w327w(0) <= wire_w_dataa_range325w(0) OR wire_w_dataa_man_not_zero_range320w(0);
	wire_w_lg_w_dataa_range331w333w(0) <= wire_w_dataa_range331w(0) OR wire_w_dataa_man_not_zero_range326w(0);
	wire_w_lg_w_dataa_range337w339w(0) <= wire_w_dataa_range337w(0) OR wire_w_dataa_man_not_zero_range332w(0);
	wire_w_lg_w_dataa_range343w345w(0) <= wire_w_dataa_range343w(0) OR wire_w_dataa_man_not_zero_range338w(0);
	wire_w_lg_w_dataa_range353w355w(0) <= wire_w_dataa_range353w(0) OR wire_w_dataa_man_not_zero_range350w(0);
	wire_w_lg_w_dataa_range359w361w(0) <= wire_w_dataa_range359w(0) OR wire_w_dataa_man_not_zero_range354w(0);
	wire_w_lg_w_dataa_range365w367w(0) <= wire_w_dataa_range365w(0) OR wire_w_dataa_man_not_zero_range360w(0);
	wire_w_lg_w_dataa_range205w207w(0) <= wire_w_dataa_range205w(0) OR wire_w_dataa_man_not_zero_range200w(0);
	wire_w_lg_w_dataa_range371w373w(0) <= wire_w_dataa_range371w(0) OR wire_w_dataa_man_not_zero_range366w(0);
	wire_w_lg_w_dataa_range377w379w(0) <= wire_w_dataa_range377w(0) OR wire_w_dataa_man_not_zero_range372w(0);
	wire_w_lg_w_dataa_range383w385w(0) <= wire_w_dataa_range383w(0) OR wire_w_dataa_man_not_zero_range378w(0);
	wire_w_lg_w_dataa_range389w391w(0) <= wire_w_dataa_range389w(0) OR wire_w_dataa_man_not_zero_range384w(0);
	wire_w_lg_w_dataa_range395w397w(0) <= wire_w_dataa_range395w(0) OR wire_w_dataa_man_not_zero_range390w(0);
	wire_w_lg_w_dataa_range401w403w(0) <= wire_w_dataa_range401w(0) OR wire_w_dataa_man_not_zero_range396w(0);
	wire_w_lg_w_dataa_range407w409w(0) <= wire_w_dataa_range407w(0) OR wire_w_dataa_man_not_zero_range402w(0);
	wire_w_lg_w_dataa_range413w415w(0) <= wire_w_dataa_range413w(0) OR wire_w_dataa_man_not_zero_range408w(0);
	wire_w_lg_w_dataa_range419w421w(0) <= wire_w_dataa_range419w(0) OR wire_w_dataa_man_not_zero_range414w(0);
	wire_w_lg_w_dataa_range425w427w(0) <= wire_w_dataa_range425w(0) OR wire_w_dataa_man_not_zero_range420w(0);
	wire_w_lg_w_dataa_range211w213w(0) <= wire_w_dataa_range211w(0) OR wire_w_dataa_man_not_zero_range206w(0);
	wire_w_lg_w_dataa_range431w433w(0) <= wire_w_dataa_range431w(0) OR wire_w_dataa_man_not_zero_range426w(0);
	wire_w_lg_w_dataa_range437w439w(0) <= wire_w_dataa_range437w(0) OR wire_w_dataa_man_not_zero_range432w(0);
	wire_w_lg_w_dataa_range443w445w(0) <= wire_w_dataa_range443w(0) OR wire_w_dataa_man_not_zero_range438w(0);
	wire_w_lg_w_dataa_range449w451w(0) <= wire_w_dataa_range449w(0) OR wire_w_dataa_man_not_zero_range444w(0);
	wire_w_lg_w_dataa_range455w457w(0) <= wire_w_dataa_range455w(0) OR wire_w_dataa_man_not_zero_range450w(0);
	wire_w_lg_w_dataa_range461w463w(0) <= wire_w_dataa_range461w(0) OR wire_w_dataa_man_not_zero_range456w(0);
	wire_w_lg_w_dataa_range467w469w(0) <= wire_w_dataa_range467w(0) OR wire_w_dataa_man_not_zero_range462w(0);
	wire_w_lg_w_dataa_range473w475w(0) <= wire_w_dataa_range473w(0) OR wire_w_dataa_man_not_zero_range468w(0);
	wire_w_lg_w_dataa_range479w481w(0) <= wire_w_dataa_range479w(0) OR wire_w_dataa_man_not_zero_range474w(0);
	wire_w_lg_w_dataa_range485w487w(0) <= wire_w_dataa_range485w(0) OR wire_w_dataa_man_not_zero_range480w(0);
	wire_w_lg_w_dataa_range217w219w(0) <= wire_w_dataa_range217w(0) OR wire_w_dataa_man_not_zero_range212w(0);
	wire_w_lg_w_dataa_range491w493w(0) <= wire_w_dataa_range491w(0) OR wire_w_dataa_man_not_zero_range486w(0);
	wire_w_lg_w_dataa_range497w499w(0) <= wire_w_dataa_range497w(0) OR wire_w_dataa_man_not_zero_range492w(0);
	wire_w_lg_w_dataa_range93w95w(0) <= wire_w_dataa_range93w(0) OR wire_w_dataa_exp_not_zero_range84w(0);
	wire_w_lg_w_dataa_range103w105w(0) <= wire_w_dataa_range103w(0) OR wire_w_dataa_exp_not_zero_range94w(0);
	wire_w_lg_w_dataa_range113w115w(0) <= wire_w_dataa_range113w(0) OR wire_w_dataa_exp_not_zero_range104w(0);
	wire_w_lg_w_dataa_range123w125w(0) <= wire_w_dataa_range123w(0) OR wire_w_dataa_exp_not_zero_range114w(0);
	wire_w_lg_w_dataa_range133w135w(0) <= wire_w_dataa_range133w(0) OR wire_w_dataa_exp_not_zero_range124w(0);
	wire_w_lg_w_dataa_range143w145w(0) <= wire_w_dataa_range143w(0) OR wire_w_dataa_exp_not_zero_range134w(0);
	wire_w_lg_w_dataa_range153w155w(0) <= wire_w_dataa_range153w(0) OR wire_w_dataa_exp_not_zero_range144w(0);
	wire_w_lg_w_dataa_range223w225w(0) <= wire_w_dataa_range223w(0) OR wire_w_dataa_man_not_zero_range218w(0);
	wire_w_lg_w_dataa_range163w165w(0) <= wire_w_dataa_range163w(0) OR wire_w_dataa_exp_not_zero_range154w(0);
	wire_w_lg_w_dataa_range173w175w(0) <= wire_w_dataa_range173w(0) OR wire_w_dataa_exp_not_zero_range164w(0);
	wire_w_lg_w_dataa_range183w185w(0) <= wire_w_dataa_range183w(0) OR wire_w_dataa_exp_not_zero_range174w(0);
	wire_w_lg_w_dataa_range229w231w(0) <= wire_w_dataa_range229w(0) OR wire_w_dataa_man_not_zero_range224w(0);
	wire_w_lg_w_dataa_range235w237w(0) <= wire_w_dataa_range235w(0) OR wire_w_dataa_man_not_zero_range230w(0);
	wire_w_lg_w_dataa_range241w243w(0) <= wire_w_dataa_range241w(0) OR wire_w_dataa_man_not_zero_range236w(0);
	wire_w_lg_w_dataa_range247w249w(0) <= wire_w_dataa_range247w(0) OR wire_w_dataa_man_not_zero_range242w(0);
	wire_w_lg_w_datab_range256w258w(0) <= wire_w_datab_range256w(0) OR wire_w_datab_man_not_zero_range251w(0);
	wire_w_lg_w_datab_range262w264w(0) <= wire_w_datab_range262w(0) OR wire_w_datab_man_not_zero_range257w(0);
	wire_w_lg_w_datab_range268w270w(0) <= wire_w_datab_range268w(0) OR wire_w_datab_man_not_zero_range263w(0);
	wire_w_lg_w_datab_range274w276w(0) <= wire_w_datab_range274w(0) OR wire_w_datab_man_not_zero_range269w(0);
	wire_w_lg_w_datab_range280w282w(0) <= wire_w_datab_range280w(0) OR wire_w_datab_man_not_zero_range275w(0);
	wire_w_lg_w_datab_range286w288w(0) <= wire_w_datab_range286w(0) OR wire_w_datab_man_not_zero_range281w(0);
	wire_w_lg_w_datab_range292w294w(0) <= wire_w_datab_range292w(0) OR wire_w_datab_man_not_zero_range287w(0);
	wire_w_lg_w_datab_range298w300w(0) <= wire_w_datab_range298w(0) OR wire_w_datab_man_not_zero_range293w(0);
	wire_w_lg_w_datab_range304w306w(0) <= wire_w_datab_range304w(0) OR wire_w_datab_man_not_zero_range299w(0);
	wire_w_lg_w_datab_range310w312w(0) <= wire_w_datab_range310w(0) OR wire_w_datab_man_not_zero_range305w(0);
	wire_w_lg_w_datab_range202w204w(0) <= wire_w_datab_range202w(0) OR wire_w_datab_man_not_zero_range197w(0);
	wire_w_lg_w_datab_range316w318w(0) <= wire_w_datab_range316w(0) OR wire_w_datab_man_not_zero_range311w(0);
	wire_w_lg_w_datab_range322w324w(0) <= wire_w_datab_range322w(0) OR wire_w_datab_man_not_zero_range317w(0);
	wire_w_lg_w_datab_range328w330w(0) <= wire_w_datab_range328w(0) OR wire_w_datab_man_not_zero_range323w(0);
	wire_w_lg_w_datab_range334w336w(0) <= wire_w_datab_range334w(0) OR wire_w_datab_man_not_zero_range329w(0);
	wire_w_lg_w_datab_range340w342w(0) <= wire_w_datab_range340w(0) OR wire_w_datab_man_not_zero_range335w(0);
	wire_w_lg_w_datab_range346w348w(0) <= wire_w_datab_range346w(0) OR wire_w_datab_man_not_zero_range341w(0);
	wire_w_lg_w_datab_range356w358w(0) <= wire_w_datab_range356w(0) OR wire_w_datab_man_not_zero_range352w(0);
	wire_w_lg_w_datab_range362w364w(0) <= wire_w_datab_range362w(0) OR wire_w_datab_man_not_zero_range357w(0);
	wire_w_lg_w_datab_range368w370w(0) <= wire_w_datab_range368w(0) OR wire_w_datab_man_not_zero_range363w(0);
	wire_w_lg_w_datab_range208w210w(0) <= wire_w_datab_range208w(0) OR wire_w_datab_man_not_zero_range203w(0);
	wire_w_lg_w_datab_range374w376w(0) <= wire_w_datab_range374w(0) OR wire_w_datab_man_not_zero_range369w(0);
	wire_w_lg_w_datab_range380w382w(0) <= wire_w_datab_range380w(0) OR wire_w_datab_man_not_zero_range375w(0);
	wire_w_lg_w_datab_range386w388w(0) <= wire_w_datab_range386w(0) OR wire_w_datab_man_not_zero_range381w(0);
	wire_w_lg_w_datab_range392w394w(0) <= wire_w_datab_range392w(0) OR wire_w_datab_man_not_zero_range387w(0);
	wire_w_lg_w_datab_range398w400w(0) <= wire_w_datab_range398w(0) OR wire_w_datab_man_not_zero_range393w(0);
	wire_w_lg_w_datab_range404w406w(0) <= wire_w_datab_range404w(0) OR wire_w_datab_man_not_zero_range399w(0);
	wire_w_lg_w_datab_range410w412w(0) <= wire_w_datab_range410w(0) OR wire_w_datab_man_not_zero_range405w(0);
	wire_w_lg_w_datab_range416w418w(0) <= wire_w_datab_range416w(0) OR wire_w_datab_man_not_zero_range411w(0);
	wire_w_lg_w_datab_range422w424w(0) <= wire_w_datab_range422w(0) OR wire_w_datab_man_not_zero_range417w(0);
	wire_w_lg_w_datab_range428w430w(0) <= wire_w_datab_range428w(0) OR wire_w_datab_man_not_zero_range423w(0);
	wire_w_lg_w_datab_range214w216w(0) <= wire_w_datab_range214w(0) OR wire_w_datab_man_not_zero_range209w(0);
	wire_w_lg_w_datab_range434w436w(0) <= wire_w_datab_range434w(0) OR wire_w_datab_man_not_zero_range429w(0);
	wire_w_lg_w_datab_range440w442w(0) <= wire_w_datab_range440w(0) OR wire_w_datab_man_not_zero_range435w(0);
	wire_w_lg_w_datab_range446w448w(0) <= wire_w_datab_range446w(0) OR wire_w_datab_man_not_zero_range441w(0);
	wire_w_lg_w_datab_range452w454w(0) <= wire_w_datab_range452w(0) OR wire_w_datab_man_not_zero_range447w(0);
	wire_w_lg_w_datab_range458w460w(0) <= wire_w_datab_range458w(0) OR wire_w_datab_man_not_zero_range453w(0);
	wire_w_lg_w_datab_range464w466w(0) <= wire_w_datab_range464w(0) OR wire_w_datab_man_not_zero_range459w(0);
	wire_w_lg_w_datab_range470w472w(0) <= wire_w_datab_range470w(0) OR wire_w_datab_man_not_zero_range465w(0);
	wire_w_lg_w_datab_range476w478w(0) <= wire_w_datab_range476w(0) OR wire_w_datab_man_not_zero_range471w(0);
	wire_w_lg_w_datab_range482w484w(0) <= wire_w_datab_range482w(0) OR wire_w_datab_man_not_zero_range477w(0);
	wire_w_lg_w_datab_range488w490w(0) <= wire_w_datab_range488w(0) OR wire_w_datab_man_not_zero_range483w(0);
	wire_w_lg_w_datab_range220w222w(0) <= wire_w_datab_range220w(0) OR wire_w_datab_man_not_zero_range215w(0);
	wire_w_lg_w_datab_range494w496w(0) <= wire_w_datab_range494w(0) OR wire_w_datab_man_not_zero_range489w(0);
	wire_w_lg_w_datab_range500w502w(0) <= wire_w_datab_range500w(0) OR wire_w_datab_man_not_zero_range495w(0);
	wire_w_lg_w_datab_range96w98w(0) <= wire_w_datab_range96w(0) OR wire_w_datab_exp_not_zero_range87w(0);
	wire_w_lg_w_datab_range106w108w(0) <= wire_w_datab_range106w(0) OR wire_w_datab_exp_not_zero_range97w(0);
	wire_w_lg_w_datab_range116w118w(0) <= wire_w_datab_range116w(0) OR wire_w_datab_exp_not_zero_range107w(0);
	wire_w_lg_w_datab_range126w128w(0) <= wire_w_datab_range126w(0) OR wire_w_datab_exp_not_zero_range117w(0);
	wire_w_lg_w_datab_range136w138w(0) <= wire_w_datab_range136w(0) OR wire_w_datab_exp_not_zero_range127w(0);
	wire_w_lg_w_datab_range146w148w(0) <= wire_w_datab_range146w(0) OR wire_w_datab_exp_not_zero_range137w(0);
	wire_w_lg_w_datab_range156w158w(0) <= wire_w_datab_range156w(0) OR wire_w_datab_exp_not_zero_range147w(0);
	wire_w_lg_w_datab_range226w228w(0) <= wire_w_datab_range226w(0) OR wire_w_datab_man_not_zero_range221w(0);
	wire_w_lg_w_datab_range166w168w(0) <= wire_w_datab_range166w(0) OR wire_w_datab_exp_not_zero_range157w(0);
	wire_w_lg_w_datab_range176w178w(0) <= wire_w_datab_range176w(0) OR wire_w_datab_exp_not_zero_range167w(0);
	wire_w_lg_w_datab_range186w188w(0) <= wire_w_datab_range186w(0) OR wire_w_datab_exp_not_zero_range177w(0);
	wire_w_lg_w_datab_range232w234w(0) <= wire_w_datab_range232w(0) OR wire_w_datab_man_not_zero_range227w(0);
	wire_w_lg_w_datab_range238w240w(0) <= wire_w_datab_range238w(0) OR wire_w_datab_man_not_zero_range233w(0);
	wire_w_lg_w_datab_range244w246w(0) <= wire_w_datab_range244w(0) OR wire_w_datab_man_not_zero_range239w(0);
	wire_w_lg_w_datab_range250w252w(0) <= wire_w_datab_range250w(0) OR wire_w_datab_man_not_zero_range245w(0);
	wire_w_lg_w_result_exp_not_zero_range745w748w(0) <= wire_w_result_exp_not_zero_range745w(0) OR wire_exp_adj_adder_w_result_range708w(0);
	wire_w_lg_w_result_exp_not_zero_range765w768w(0) <= wire_w_result_exp_not_zero_range765w(0) OR wire_exp_adj_adder_w_result_range738w(0);
	wire_w_lg_w_result_exp_not_zero_range747w750w(0) <= wire_w_result_exp_not_zero_range747w(0) OR wire_exp_adj_adder_w_result_range711w(0);
	wire_w_lg_w_result_exp_not_zero_range749w752w(0) <= wire_w_result_exp_not_zero_range749w(0) OR wire_exp_adj_adder_w_result_range714w(0);
	wire_w_lg_w_result_exp_not_zero_range751w754w(0) <= wire_w_result_exp_not_zero_range751w(0) OR wire_exp_adj_adder_w_result_range717w(0);
	wire_w_lg_w_result_exp_not_zero_range753w756w(0) <= wire_w_result_exp_not_zero_range753w(0) OR wire_exp_adj_adder_w_result_range720w(0);
	wire_w_lg_w_result_exp_not_zero_range755w758w(0) <= wire_w_result_exp_not_zero_range755w(0) OR wire_exp_adj_adder_w_result_range723w(0);
	wire_w_lg_w_result_exp_not_zero_range757w760w(0) <= wire_w_result_exp_not_zero_range757w(0) OR wire_exp_adj_adder_w_result_range726w(0);
	wire_w_lg_w_result_exp_not_zero_range759w762w(0) <= wire_w_result_exp_not_zero_range759w(0) OR wire_exp_adj_adder_w_result_range729w(0);
	wire_w_lg_w_result_exp_not_zero_range761w764w(0) <= wire_w_result_exp_not_zero_range761w(0) OR wire_exp_adj_adder_w_result_range732w(0);
	wire_w_lg_w_result_exp_not_zero_range763w766w(0) <= wire_w_result_exp_not_zero_range763w(0) OR wire_exp_adj_adder_w_result_range735w(0);
	wire_w_lg_w_sticky_bit_range522w526w(0) <= wire_w_sticky_bit_range522w(0) OR wire_man_product2_mult_w_result_range524w(0);
	wire_w_lg_w_sticky_bit_range552w556w(0) <= wire_w_sticky_bit_range552w(0) OR wire_man_product2_mult_w_result_range554w(0);
	wire_w_lg_w_sticky_bit_range555w559w(0) <= wire_w_sticky_bit_range555w(0) OR wire_man_product2_mult_w_result_range557w(0);
	wire_w_lg_w_sticky_bit_range558w562w(0) <= wire_w_sticky_bit_range558w(0) OR wire_man_product2_mult_w_result_range560w(0);
	wire_w_lg_w_sticky_bit_range561w565w(0) <= wire_w_sticky_bit_range561w(0) OR wire_man_product2_mult_w_result_range563w(0);
	wire_w_lg_w_sticky_bit_range564w568w(0) <= wire_w_sticky_bit_range564w(0) OR wire_man_product2_mult_w_result_range566w(0);
	wire_w_lg_w_sticky_bit_range567w571w(0) <= wire_w_sticky_bit_range567w(0) OR wire_man_product2_mult_w_result_range569w(0);
	wire_w_lg_w_sticky_bit_range570w574w(0) <= wire_w_sticky_bit_range570w(0) OR wire_man_product2_mult_w_result_range572w(0);
	wire_w_lg_w_sticky_bit_range573w577w(0) <= wire_w_sticky_bit_range573w(0) OR wire_man_product2_mult_w_result_range575w(0);
	wire_w_lg_w_sticky_bit_range576w580w(0) <= wire_w_sticky_bit_range576w(0) OR wire_man_product2_mult_w_result_range578w(0);
	wire_w_lg_w_sticky_bit_range579w583w(0) <= wire_w_sticky_bit_range579w(0) OR wire_man_product2_mult_w_result_range581w(0);
	wire_w_lg_w_sticky_bit_range525w529w(0) <= wire_w_sticky_bit_range525w(0) OR wire_man_product2_mult_w_result_range527w(0);
	wire_w_lg_w_sticky_bit_range582w586w(0) <= wire_w_sticky_bit_range582w(0) OR wire_man_product2_mult_w_result_range584w(0);
	wire_w_lg_w_sticky_bit_range585w589w(0) <= wire_w_sticky_bit_range585w(0) OR wire_man_product2_mult_w_result_range587w(0);
	wire_w_lg_w_sticky_bit_range588w592w(0) <= wire_w_sticky_bit_range588w(0) OR wire_man_product2_mult_w_result_range590w(0);
	wire_w_lg_w_sticky_bit_range591w595w(0) <= wire_w_sticky_bit_range591w(0) OR wire_man_product2_mult_w_result_range593w(0);
	wire_w_lg_w_sticky_bit_range594w598w(0) <= wire_w_sticky_bit_range594w(0) OR wire_man_product2_mult_w_result_range596w(0);
	wire_w_lg_w_sticky_bit_range597w601w(0) <= wire_w_sticky_bit_range597w(0) OR wire_man_product2_mult_w_result_range599w(0);
	wire_w_lg_w_sticky_bit_range600w604w(0) <= wire_w_sticky_bit_range600w(0) OR wire_man_product2_mult_w_result_range602w(0);
	wire_w_lg_w_sticky_bit_range603w607w(0) <= wire_w_sticky_bit_range603w(0) OR wire_man_product2_mult_w_result_range605w(0);
	wire_w_lg_w_sticky_bit_range606w610w(0) <= wire_w_sticky_bit_range606w(0) OR wire_man_product2_mult_w_result_range608w(0);
	wire_w_lg_w_sticky_bit_range609w613w(0) <= wire_w_sticky_bit_range609w(0) OR wire_man_product2_mult_w_result_range611w(0);
	wire_w_lg_w_sticky_bit_range528w532w(0) <= wire_w_sticky_bit_range528w(0) OR wire_man_product2_mult_w_result_range530w(0);
	wire_w_lg_w_sticky_bit_range612w616w(0) <= wire_w_sticky_bit_range612w(0) OR wire_man_product2_mult_w_result_range614w(0);
	wire_w_lg_w_sticky_bit_range615w619w(0) <= wire_w_sticky_bit_range615w(0) OR wire_man_product2_mult_w_result_range617w(0);
	wire_w_lg_w_sticky_bit_range618w622w(0) <= wire_w_sticky_bit_range618w(0) OR wire_man_product2_mult_w_result_range620w(0);
	wire_w_lg_w_sticky_bit_range621w625w(0) <= wire_w_sticky_bit_range621w(0) OR wire_man_product2_mult_w_result_range623w(0);
	wire_w_lg_w_sticky_bit_range624w628w(0) <= wire_w_sticky_bit_range624w(0) OR wire_man_product2_mult_w_result_range626w(0);
	wire_w_lg_w_sticky_bit_range627w631w(0) <= wire_w_sticky_bit_range627w(0) OR wire_man_product2_mult_w_result_range629w(0);
	wire_w_lg_w_sticky_bit_range630w634w(0) <= wire_w_sticky_bit_range630w(0) OR wire_man_product2_mult_w_result_range632w(0);
	wire_w_lg_w_sticky_bit_range633w637w(0) <= wire_w_sticky_bit_range633w(0) OR wire_man_product2_mult_w_result_range635w(0);
	wire_w_lg_w_sticky_bit_range636w640w(0) <= wire_w_sticky_bit_range636w(0) OR wire_man_product2_mult_w_result_range638w(0);
	wire_w_lg_w_sticky_bit_range639w643w(0) <= wire_w_sticky_bit_range639w(0) OR wire_man_product2_mult_w_result_range641w(0);
	wire_w_lg_w_sticky_bit_range531w535w(0) <= wire_w_sticky_bit_range531w(0) OR wire_man_product2_mult_w_result_range533w(0);
	wire_w_lg_w_sticky_bit_range642w646w(0) <= wire_w_sticky_bit_range642w(0) OR wire_man_product2_mult_w_result_range644w(0);
	wire_w_lg_w_sticky_bit_range645w649w(0) <= wire_w_sticky_bit_range645w(0) OR wire_man_product2_mult_w_result_range647w(0);
	wire_w_lg_w_sticky_bit_range648w652w(0) <= wire_w_sticky_bit_range648w(0) OR wire_man_product2_mult_w_result_range650w(0);
	wire_w_lg_w_sticky_bit_range651w655w(0) <= wire_w_sticky_bit_range651w(0) OR wire_man_product2_mult_w_result_range653w(0);
	wire_w_lg_w_sticky_bit_range654w658w(0) <= wire_w_sticky_bit_range654w(0) OR wire_man_product2_mult_w_result_range656w(0);
	wire_w_lg_w_sticky_bit_range657w661w(0) <= wire_w_sticky_bit_range657w(0) OR wire_man_product2_mult_w_result_range659w(0);
	wire_w_lg_w_sticky_bit_range660w664w(0) <= wire_w_sticky_bit_range660w(0) OR wire_man_product2_mult_w_result_range662w(0);
	wire_w_lg_w_sticky_bit_range663w667w(0) <= wire_w_sticky_bit_range663w(0) OR wire_man_product2_mult_w_result_range665w(0);
	wire_w_lg_w_sticky_bit_range666w670w(0) <= wire_w_sticky_bit_range666w(0) OR wire_man_product2_mult_w_result_range668w(0);
	wire_w_lg_w_sticky_bit_range669w673w(0) <= wire_w_sticky_bit_range669w(0) OR wire_man_product2_mult_w_result_range671w(0);
	wire_w_lg_w_sticky_bit_range534w538w(0) <= wire_w_sticky_bit_range534w(0) OR wire_man_product2_mult_w_result_range536w(0);
	wire_w_lg_w_sticky_bit_range672w677w(0) <= wire_w_sticky_bit_range672w(0) OR wire_man_product2_mult_w_lg_w_result_range514w676w(0);
	wire_w_lg_w_sticky_bit_range537w541w(0) <= wire_w_sticky_bit_range537w(0) OR wire_man_product2_mult_w_result_range539w(0);
	wire_w_lg_w_sticky_bit_range540w544w(0) <= wire_w_sticky_bit_range540w(0) OR wire_man_product2_mult_w_result_range542w(0);
	wire_w_lg_w_sticky_bit_range543w547w(0) <= wire_w_sticky_bit_range543w(0) OR wire_man_product2_mult_w_result_range545w(0);
	wire_w_lg_w_sticky_bit_range546w550w(0) <= wire_w_sticky_bit_range546w(0) OR wire_man_product2_mult_w_result_range548w(0);
	wire_w_lg_w_sticky_bit_range549w553w(0) <= wire_w_sticky_bit_range549w(0) OR wire_man_product2_mult_w_result_range551w(0);
	aclr <= '0';
	bias <= ( "0" & "0" & "0" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1");
	clk_en <= '1';
	dataa_exp_all_one <= ( wire_w_lg_w_dataa_range183w190w & wire_w_lg_w_dataa_range173w180w & wire_w_lg_w_dataa_range163w170w & wire_w_lg_w_dataa_range153w160w & wire_w_lg_w_dataa_range143w150w & wire_w_lg_w_dataa_range133w140w & wire_w_lg_w_dataa_range123w130w & wire_w_lg_w_dataa_range113w120w & wire_w_lg_w_dataa_range103w110w & wire_w_lg_w_dataa_range93w100w & dataa(52));
	dataa_exp_not_zero <= ( wire_w_lg_w_dataa_range183w185w & wire_w_lg_w_dataa_range173w175w & wire_w_lg_w_dataa_range163w165w & wire_w_lg_w_dataa_range153w155w & wire_w_lg_w_dataa_range143w145w & wire_w_lg_w_dataa_range133w135w & wire_w_lg_w_dataa_range123w125w & wire_w_lg_w_dataa_range113w115w & wire_w_lg_w_dataa_range103w105w & wire_w_lg_w_dataa_range93w95w & dataa(52));
	dataa_man_not_zero <= ( wire_w_lg_w_dataa_range497w499w & wire_w_lg_w_dataa_range491w493w & wire_w_lg_w_dataa_range485w487w & wire_w_lg_w_dataa_range479w481w & wire_w_lg_w_dataa_range473w475w & wire_w_lg_w_dataa_range467w469w & wire_w_lg_w_dataa_range461w463w & wire_w_lg_w_dataa_range455w457w & wire_w_lg_w_dataa_range449w451w & wire_w_lg_w_dataa_range443w445w & wire_w_lg_w_dataa_range437w439w & wire_w_lg_w_dataa_range431w433w & wire_w_lg_w_dataa_range425w427w & wire_w_lg_w_dataa_range419w421w & wire_w_lg_w_dataa_range413w415w & wire_w_lg_w_dataa_range407w409w & wire_w_lg_w_dataa_range401w403w & wire_w_lg_w_dataa_range395w397w & wire_w_lg_w_dataa_range389w391w & wire_w_lg_w_dataa_range383w385w & wire_w_lg_w_dataa_range377w379w & wire_w_lg_w_dataa_range371w373w & wire_w_lg_w_dataa_range365w367w & wire_w_lg_w_dataa_range359w361w & wire_w_lg_w_dataa_range353w355w & dataa(26) & wire_w_lg_w_dataa_range343w345w & wire_w_lg_w_dataa_range337w339w & wire_w_lg_w_dataa_range331w333w & wire_w_lg_w_dataa_range325w327w & wire_w_lg_w_dataa_range319w321w & wire_w_lg_w_dataa_range313w315w & wire_w_lg_w_dataa_range307w309w & wire_w_lg_w_dataa_range301w303w & wire_w_lg_w_dataa_range295w297w & wire_w_lg_w_dataa_range289w291w & wire_w_lg_w_dataa_range283w285w & wire_w_lg_w_dataa_range277w279w & wire_w_lg_w_dataa_range271w273w & wire_w_lg_w_dataa_range265w267w & wire_w_lg_w_dataa_range259w261w & wire_w_lg_w_dataa_range253w255w & wire_w_lg_w_dataa_range247w249w & wire_w_lg_w_dataa_range241w243w & wire_w_lg_w_dataa_range235w237w & wire_w_lg_w_dataa_range229w231w & wire_w_lg_w_dataa_range223w225w & wire_w_lg_w_dataa_range217w219w & wire_w_lg_w_dataa_range211w213w & wire_w_lg_w_dataa_range205w207w & wire_w_lg_w_dataa_range199w201w & dataa(0));
	datab_exp_all_one <= ( wire_w_lg_w_datab_range186w192w & wire_w_lg_w_datab_range176w182w & wire_w_lg_w_datab_range166w172w & wire_w_lg_w_datab_range156w162w & wire_w_lg_w_datab_range146w152w & wire_w_lg_w_datab_range136w142w & wire_w_lg_w_datab_range126w132w & wire_w_lg_w_datab_range116w122w & wire_w_lg_w_datab_range106w112w & wire_w_lg_w_datab_range96w102w & datab(52));
	datab_exp_not_zero <= ( wire_w_lg_w_datab_range186w188w & wire_w_lg_w_datab_range176w178w & wire_w_lg_w_datab_range166w168w & wire_w_lg_w_datab_range156w158w & wire_w_lg_w_datab_range146w148w & wire_w_lg_w_datab_range136w138w & wire_w_lg_w_datab_range126w128w & wire_w_lg_w_datab_range116w118w & wire_w_lg_w_datab_range106w108w & wire_w_lg_w_datab_range96w98w & datab(52));
	datab_man_not_zero <= ( wire_w_lg_w_datab_range500w502w & wire_w_lg_w_datab_range494w496w & wire_w_lg_w_datab_range488w490w & wire_w_lg_w_datab_range482w484w & wire_w_lg_w_datab_range476w478w & wire_w_lg_w_datab_range470w472w & wire_w_lg_w_datab_range464w466w & wire_w_lg_w_datab_range458w460w & wire_w_lg_w_datab_range452w454w & wire_w_lg_w_datab_range446w448w & wire_w_lg_w_datab_range440w442w & wire_w_lg_w_datab_range434w436w & wire_w_lg_w_datab_range428w430w & wire_w_lg_w_datab_range422w424w & wire_w_lg_w_datab_range416w418w & wire_w_lg_w_datab_range410w412w & wire_w_lg_w_datab_range404w406w & wire_w_lg_w_datab_range398w400w & wire_w_lg_w_datab_range392w394w & wire_w_lg_w_datab_range386w388w & wire_w_lg_w_datab_range380w382w & wire_w_lg_w_datab_range374w376w & wire_w_lg_w_datab_range368w370w & wire_w_lg_w_datab_range362w364w & wire_w_lg_w_datab_range356w358w & datab(26) & wire_w_lg_w_datab_range346w348w & wire_w_lg_w_datab_range340w342w & wire_w_lg_w_datab_range334w336w & wire_w_lg_w_datab_range328w330w & wire_w_lg_w_datab_range322w324w & wire_w_lg_w_datab_range316w318w & wire_w_lg_w_datab_range310w312w & wire_w_lg_w_datab_range304w306w & wire_w_lg_w_datab_range298w300w & wire_w_lg_w_datab_range292w294w & wire_w_lg_w_datab_range286w288w & wire_w_lg_w_datab_range280w282w & wire_w_lg_w_datab_range274w276w & wire_w_lg_w_datab_range268w270w & wire_w_lg_w_datab_range262w264w & wire_w_lg_w_datab_range256w258w & wire_w_lg_w_datab_range250w252w & wire_w_lg_w_datab_range244w246w & wire_w_lg_w_datab_range238w240w & wire_w_lg_w_datab_range232w234w & wire_w_lg_w_datab_range226w228w & wire_w_lg_w_datab_range220w222w & wire_w_lg_w_datab_range214w216w & wire_w_lg_w_datab_range208w210w & wire_w_lg_w_datab_range202w204w & datab(0));
	exp_is_inf <= (((NOT wire_exp_adj_adder_result(12)) AND wire_exp_adj_adder_result(11)) OR ((NOT wire_exp_adj_adder_result(11)) AND result_exp_all_one(10)));
	exp_is_zero <= wire_exp_adj_adder_w_lg_w_result_range739w770w(0);
	expmod <= ( "00000000000" & wire_delay_man_product_msb_w_lg_q696w & wire_delay_man_product_msb_w_lg_q698w);
	inf_num <= ( "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1");
	lsb_bit <= man_shift_full(1);
	man_result_round <= (wire_man_round_p2_w_lg_w_q_range702w703w OR wire_man_round_p2_w_lg_w_q_range699w700w);
	man_shift_full <= (wire_man_product2_mult_w_lg_w_result_range518w519w OR wire_man_product2_mult_w_lg_w_result_range515w516w);
	overflow <= overflow_ff;
	result <= ( sign_node_ff4 & exp_result_ff(10 DOWNTO 0) & man_result_ff(51 DOWNTO 0));
	result_exp_all_one <= ( wire_w_lg_w_result_exp_all_one_range733w737w & wire_w_lg_w_result_exp_all_one_range730w734w & wire_w_lg_w_result_exp_all_one_range727w731w & wire_w_lg_w_result_exp_all_one_range724w728w & wire_w_lg_w_result_exp_all_one_range721w725w & wire_w_lg_w_result_exp_all_one_range718w722w & wire_w_lg_w_result_exp_all_one_range715w719w & wire_w_lg_w_result_exp_all_one_range712w716w & wire_w_lg_w_result_exp_all_one_range709w713w & wire_w_lg_w_result_exp_all_one_range706w710w & wire_exp_adj_adder_result(0));
	result_exp_not_zero <= ( wire_w_lg_w_result_exp_not_zero_range765w768w & wire_w_lg_w_result_exp_not_zero_range763w766w & wire_w_lg_w_result_exp_not_zero_range761w764w & wire_w_lg_w_result_exp_not_zero_range759w762w & wire_w_lg_w_result_exp_not_zero_range757w760w & wire_w_lg_w_result_exp_not_zero_range755w758w & wire_w_lg_w_result_exp_not_zero_range753w756w & wire_w_lg_w_result_exp_not_zero_range751w754w & wire_w_lg_w_result_exp_not_zero_range749w752w & wire_w_lg_w_result_exp_not_zero_range747w750w & wire_w_lg_w_result_exp_not_zero_range745w748w & wire_exp_adj_adder_result(0));
	round_bit <= man_shift_full(0);
	round_carry <= (round_dffe AND (lsb_dffe OR sticky_dffe));
	sticky_bit <= ( wire_w_lg_w_sticky_bit_range672w677w & wire_w_lg_w_sticky_bit_range669w673w & wire_w_lg_w_sticky_bit_range666w670w & wire_w_lg_w_sticky_bit_range663w667w & wire_w_lg_w_sticky_bit_range660w664w & wire_w_lg_w_sticky_bit_range657w661w & wire_w_lg_w_sticky_bit_range654w658w & wire_w_lg_w_sticky_bit_range651w655w & wire_w_lg_w_sticky_bit_range648w652w & wire_w_lg_w_sticky_bit_range645w649w & wire_w_lg_w_sticky_bit_range642w646w & wire_w_lg_w_sticky_bit_range639w643w & wire_w_lg_w_sticky_bit_range636w640w & wire_w_lg_w_sticky_bit_range633w637w & wire_w_lg_w_sticky_bit_range630w634w & wire_w_lg_w_sticky_bit_range627w631w & wire_w_lg_w_sticky_bit_range624w628w & wire_w_lg_w_sticky_bit_range621w625w & wire_w_lg_w_sticky_bit_range618w622w & wire_w_lg_w_sticky_bit_range615w619w & wire_w_lg_w_sticky_bit_range612w616w & wire_w_lg_w_sticky_bit_range609w613w & wire_w_lg_w_sticky_bit_range606w610w & wire_w_lg_w_sticky_bit_range603w607w & wire_w_lg_w_sticky_bit_range600w604w & wire_w_lg_w_sticky_bit_range597w601w & wire_w_lg_w_sticky_bit_range594w598w & wire_w_lg_w_sticky_bit_range591w595w & wire_w_lg_w_sticky_bit_range588w592w & wire_w_lg_w_sticky_bit_range585w589w & wire_w_lg_w_sticky_bit_range582w586w & wire_w_lg_w_sticky_bit_range579w583w & wire_w_lg_w_sticky_bit_range576w580w & wire_w_lg_w_sticky_bit_range573w577w & wire_w_lg_w_sticky_bit_range570w574w & wire_w_lg_w_sticky_bit_range567w571w & wire_w_lg_w_sticky_bit_range564w568w & wire_w_lg_w_sticky_bit_range561w565w & wire_w_lg_w_sticky_bit_range558w562w & wire_w_lg_w_sticky_bit_range555w559w & wire_w_lg_w_sticky_bit_range552w556w & wire_w_lg_w_sticky_bit_range549w553w & wire_w_lg_w_sticky_bit_range546w550w & wire_w_lg_w_sticky_bit_range543w547w & wire_w_lg_w_sticky_bit_range540w544w & wire_w_lg_w_sticky_bit_range537w541w & wire_w_lg_w_sticky_bit_range534w538w & wire_w_lg_w_sticky_bit_range531w535w & wire_w_lg_w_sticky_bit_range528w532w & wire_w_lg_w_sticky_bit_range525w529w & wire_w_lg_w_sticky_bit_range522w526w & wire_man_product2_mult_result(0));
	wire_w_dataa_range253w(0) <= dataa(10);
	wire_w_dataa_range259w(0) <= dataa(11);
	wire_w_dataa_range265w(0) <= dataa(12);
	wire_w_dataa_range271w(0) <= dataa(13);
	wire_w_dataa_range277w(0) <= dataa(14);
	wire_w_dataa_range283w(0) <= dataa(15);
	wire_w_dataa_range289w(0) <= dataa(16);
	wire_w_dataa_range295w(0) <= dataa(17);
	wire_w_dataa_range301w(0) <= dataa(18);
	wire_w_dataa_range307w(0) <= dataa(19);
	wire_w_dataa_range199w(0) <= dataa(1);
	wire_w_dataa_range313w(0) <= dataa(20);
	wire_w_dataa_range319w(0) <= dataa(21);
	wire_w_dataa_range325w(0) <= dataa(22);
	wire_w_dataa_range331w(0) <= dataa(23);
	wire_w_dataa_range337w(0) <= dataa(24);
	wire_w_dataa_range343w(0) <= dataa(25);
	wire_w_dataa_range353w(0) <= dataa(27);
	wire_w_dataa_range359w(0) <= dataa(28);
	wire_w_dataa_range365w(0) <= dataa(29);
	wire_w_dataa_range205w(0) <= dataa(2);
	wire_w_dataa_range371w(0) <= dataa(30);
	wire_w_dataa_range377w(0) <= dataa(31);
	wire_w_dataa_range383w(0) <= dataa(32);
	wire_w_dataa_range389w(0) <= dataa(33);
	wire_w_dataa_range395w(0) <= dataa(34);
	wire_w_dataa_range401w(0) <= dataa(35);
	wire_w_dataa_range407w(0) <= dataa(36);
	wire_w_dataa_range413w(0) <= dataa(37);
	wire_w_dataa_range419w(0) <= dataa(38);
	wire_w_dataa_range425w(0) <= dataa(39);
	wire_w_dataa_range211w(0) <= dataa(3);
	wire_w_dataa_range431w(0) <= dataa(40);
	wire_w_dataa_range437w(0) <= dataa(41);
	wire_w_dataa_range443w(0) <= dataa(42);
	wire_w_dataa_range449w(0) <= dataa(43);
	wire_w_dataa_range455w(0) <= dataa(44);
	wire_w_dataa_range461w(0) <= dataa(45);
	wire_w_dataa_range467w(0) <= dataa(46);
	wire_w_dataa_range473w(0) <= dataa(47);
	wire_w_dataa_range479w(0) <= dataa(48);
	wire_w_dataa_range485w(0) <= dataa(49);
	wire_w_dataa_range217w(0) <= dataa(4);
	wire_w_dataa_range491w(0) <= dataa(50);
	wire_w_dataa_range497w(0) <= dataa(51);
	wire_w_dataa_range93w(0) <= dataa(53);
	wire_w_dataa_range103w(0) <= dataa(54);
	wire_w_dataa_range113w(0) <= dataa(55);
	wire_w_dataa_range123w(0) <= dataa(56);
	wire_w_dataa_range133w(0) <= dataa(57);
	wire_w_dataa_range143w(0) <= dataa(58);
	wire_w_dataa_range153w(0) <= dataa(59);
	wire_w_dataa_range223w(0) <= dataa(5);
	wire_w_dataa_range163w(0) <= dataa(60);
	wire_w_dataa_range173w(0) <= dataa(61);
	wire_w_dataa_range183w(0) <= dataa(62);
	wire_w_dataa_range229w(0) <= dataa(6);
	wire_w_dataa_range235w(0) <= dataa(7);
	wire_w_dataa_range241w(0) <= dataa(8);
	wire_w_dataa_range247w(0) <= dataa(9);
	wire_w_dataa_exp_all_one_range89w(0) <= dataa_exp_all_one(0);
	wire_w_dataa_exp_all_one_range99w(0) <= dataa_exp_all_one(1);
	wire_w_dataa_exp_all_one_range109w(0) <= dataa_exp_all_one(2);
	wire_w_dataa_exp_all_one_range119w(0) <= dataa_exp_all_one(3);
	wire_w_dataa_exp_all_one_range129w(0) <= dataa_exp_all_one(4);
	wire_w_dataa_exp_all_one_range139w(0) <= dataa_exp_all_one(5);
	wire_w_dataa_exp_all_one_range149w(0) <= dataa_exp_all_one(6);
	wire_w_dataa_exp_all_one_range159w(0) <= dataa_exp_all_one(7);
	wire_w_dataa_exp_all_one_range169w(0) <= dataa_exp_all_one(8);
	wire_w_dataa_exp_all_one_range179w(0) <= dataa_exp_all_one(9);
	wire_w_dataa_exp_not_zero_range84w(0) <= dataa_exp_not_zero(0);
	wire_w_dataa_exp_not_zero_range94w(0) <= dataa_exp_not_zero(1);
	wire_w_dataa_exp_not_zero_range104w(0) <= dataa_exp_not_zero(2);
	wire_w_dataa_exp_not_zero_range114w(0) <= dataa_exp_not_zero(3);
	wire_w_dataa_exp_not_zero_range124w(0) <= dataa_exp_not_zero(4);
	wire_w_dataa_exp_not_zero_range134w(0) <= dataa_exp_not_zero(5);
	wire_w_dataa_exp_not_zero_range144w(0) <= dataa_exp_not_zero(6);
	wire_w_dataa_exp_not_zero_range154w(0) <= dataa_exp_not_zero(7);
	wire_w_dataa_exp_not_zero_range164w(0) <= dataa_exp_not_zero(8);
	wire_w_dataa_exp_not_zero_range174w(0) <= dataa_exp_not_zero(9);
	wire_w_dataa_man_not_zero_range194w(0) <= dataa_man_not_zero(0);
	wire_w_dataa_man_not_zero_range254w(0) <= dataa_man_not_zero(10);
	wire_w_dataa_man_not_zero_range260w(0) <= dataa_man_not_zero(11);
	wire_w_dataa_man_not_zero_range266w(0) <= dataa_man_not_zero(12);
	wire_w_dataa_man_not_zero_range272w(0) <= dataa_man_not_zero(13);
	wire_w_dataa_man_not_zero_range278w(0) <= dataa_man_not_zero(14);
	wire_w_dataa_man_not_zero_range284w(0) <= dataa_man_not_zero(15);
	wire_w_dataa_man_not_zero_range290w(0) <= dataa_man_not_zero(16);
	wire_w_dataa_man_not_zero_range296w(0) <= dataa_man_not_zero(17);
	wire_w_dataa_man_not_zero_range302w(0) <= dataa_man_not_zero(18);
	wire_w_dataa_man_not_zero_range308w(0) <= dataa_man_not_zero(19);
	wire_w_dataa_man_not_zero_range200w(0) <= dataa_man_not_zero(1);
	wire_w_dataa_man_not_zero_range314w(0) <= dataa_man_not_zero(20);
	wire_w_dataa_man_not_zero_range320w(0) <= dataa_man_not_zero(21);
	wire_w_dataa_man_not_zero_range326w(0) <= dataa_man_not_zero(22);
	wire_w_dataa_man_not_zero_range332w(0) <= dataa_man_not_zero(23);
	wire_w_dataa_man_not_zero_range338w(0) <= dataa_man_not_zero(24);
	wire_w_dataa_man_not_zero_range350w(0) <= dataa_man_not_zero(26);
	wire_w_dataa_man_not_zero_range354w(0) <= dataa_man_not_zero(27);
	wire_w_dataa_man_not_zero_range360w(0) <= dataa_man_not_zero(28);
	wire_w_dataa_man_not_zero_range366w(0) <= dataa_man_not_zero(29);
	wire_w_dataa_man_not_zero_range206w(0) <= dataa_man_not_zero(2);
	wire_w_dataa_man_not_zero_range372w(0) <= dataa_man_not_zero(30);
	wire_w_dataa_man_not_zero_range378w(0) <= dataa_man_not_zero(31);
	wire_w_dataa_man_not_zero_range384w(0) <= dataa_man_not_zero(32);
	wire_w_dataa_man_not_zero_range390w(0) <= dataa_man_not_zero(33);
	wire_w_dataa_man_not_zero_range396w(0) <= dataa_man_not_zero(34);
	wire_w_dataa_man_not_zero_range402w(0) <= dataa_man_not_zero(35);
	wire_w_dataa_man_not_zero_range408w(0) <= dataa_man_not_zero(36);
	wire_w_dataa_man_not_zero_range414w(0) <= dataa_man_not_zero(37);
	wire_w_dataa_man_not_zero_range420w(0) <= dataa_man_not_zero(38);
	wire_w_dataa_man_not_zero_range426w(0) <= dataa_man_not_zero(39);
	wire_w_dataa_man_not_zero_range212w(0) <= dataa_man_not_zero(3);
	wire_w_dataa_man_not_zero_range432w(0) <= dataa_man_not_zero(40);
	wire_w_dataa_man_not_zero_range438w(0) <= dataa_man_not_zero(41);
	wire_w_dataa_man_not_zero_range444w(0) <= dataa_man_not_zero(42);
	wire_w_dataa_man_not_zero_range450w(0) <= dataa_man_not_zero(43);
	wire_w_dataa_man_not_zero_range456w(0) <= dataa_man_not_zero(44);
	wire_w_dataa_man_not_zero_range462w(0) <= dataa_man_not_zero(45);
	wire_w_dataa_man_not_zero_range468w(0) <= dataa_man_not_zero(46);
	wire_w_dataa_man_not_zero_range474w(0) <= dataa_man_not_zero(47);
	wire_w_dataa_man_not_zero_range480w(0) <= dataa_man_not_zero(48);
	wire_w_dataa_man_not_zero_range486w(0) <= dataa_man_not_zero(49);
	wire_w_dataa_man_not_zero_range218w(0) <= dataa_man_not_zero(4);
	wire_w_dataa_man_not_zero_range492w(0) <= dataa_man_not_zero(50);
	wire_w_dataa_man_not_zero_range224w(0) <= dataa_man_not_zero(5);
	wire_w_dataa_man_not_zero_range230w(0) <= dataa_man_not_zero(6);
	wire_w_dataa_man_not_zero_range236w(0) <= dataa_man_not_zero(7);
	wire_w_dataa_man_not_zero_range242w(0) <= dataa_man_not_zero(8);
	wire_w_dataa_man_not_zero_range248w(0) <= dataa_man_not_zero(9);
	wire_w_datab_range256w(0) <= datab(10);
	wire_w_datab_range262w(0) <= datab(11);
	wire_w_datab_range268w(0) <= datab(12);
	wire_w_datab_range274w(0) <= datab(13);
	wire_w_datab_range280w(0) <= datab(14);
	wire_w_datab_range286w(0) <= datab(15);
	wire_w_datab_range292w(0) <= datab(16);
	wire_w_datab_range298w(0) <= datab(17);
	wire_w_datab_range304w(0) <= datab(18);
	wire_w_datab_range310w(0) <= datab(19);
	wire_w_datab_range202w(0) <= datab(1);
	wire_w_datab_range316w(0) <= datab(20);
	wire_w_datab_range322w(0) <= datab(21);
	wire_w_datab_range328w(0) <= datab(22);
	wire_w_datab_range334w(0) <= datab(23);
	wire_w_datab_range340w(0) <= datab(24);
	wire_w_datab_range346w(0) <= datab(25);
	wire_w_datab_range356w(0) <= datab(27);
	wire_w_datab_range362w(0) <= datab(28);
	wire_w_datab_range368w(0) <= datab(29);
	wire_w_datab_range208w(0) <= datab(2);
	wire_w_datab_range374w(0) <= datab(30);
	wire_w_datab_range380w(0) <= datab(31);
	wire_w_datab_range386w(0) <= datab(32);
	wire_w_datab_range392w(0) <= datab(33);
	wire_w_datab_range398w(0) <= datab(34);
	wire_w_datab_range404w(0) <= datab(35);
	wire_w_datab_range410w(0) <= datab(36);
	wire_w_datab_range416w(0) <= datab(37);
	wire_w_datab_range422w(0) <= datab(38);
	wire_w_datab_range428w(0) <= datab(39);
	wire_w_datab_range214w(0) <= datab(3);
	wire_w_datab_range434w(0) <= datab(40);
	wire_w_datab_range440w(0) <= datab(41);
	wire_w_datab_range446w(0) <= datab(42);
	wire_w_datab_range452w(0) <= datab(43);
	wire_w_datab_range458w(0) <= datab(44);
	wire_w_datab_range464w(0) <= datab(45);
	wire_w_datab_range470w(0) <= datab(46);
	wire_w_datab_range476w(0) <= datab(47);
	wire_w_datab_range482w(0) <= datab(48);
	wire_w_datab_range488w(0) <= datab(49);
	wire_w_datab_range220w(0) <= datab(4);
	wire_w_datab_range494w(0) <= datab(50);
	wire_w_datab_range500w(0) <= datab(51);
	wire_w_datab_range96w(0) <= datab(53);
	wire_w_datab_range106w(0) <= datab(54);
	wire_w_datab_range116w(0) <= datab(55);
	wire_w_datab_range126w(0) <= datab(56);
	wire_w_datab_range136w(0) <= datab(57);
	wire_w_datab_range146w(0) <= datab(58);
	wire_w_datab_range156w(0) <= datab(59);
	wire_w_datab_range226w(0) <= datab(5);
	wire_w_datab_range166w(0) <= datab(60);
	wire_w_datab_range176w(0) <= datab(61);
	wire_w_datab_range186w(0) <= datab(62);
	wire_w_datab_range232w(0) <= datab(6);
	wire_w_datab_range238w(0) <= datab(7);
	wire_w_datab_range244w(0) <= datab(8);
	wire_w_datab_range250w(0) <= datab(9);
	wire_w_datab_exp_all_one_range91w(0) <= datab_exp_all_one(0);
	wire_w_datab_exp_all_one_range101w(0) <= datab_exp_all_one(1);
	wire_w_datab_exp_all_one_range111w(0) <= datab_exp_all_one(2);
	wire_w_datab_exp_all_one_range121w(0) <= datab_exp_all_one(3);
	wire_w_datab_exp_all_one_range131w(0) <= datab_exp_all_one(4);
	wire_w_datab_exp_all_one_range141w(0) <= datab_exp_all_one(5);
	wire_w_datab_exp_all_one_range151w(0) <= datab_exp_all_one(6);
	wire_w_datab_exp_all_one_range161w(0) <= datab_exp_all_one(7);
	wire_w_datab_exp_all_one_range171w(0) <= datab_exp_all_one(8);
	wire_w_datab_exp_all_one_range181w(0) <= datab_exp_all_one(9);
	wire_w_datab_exp_not_zero_range87w(0) <= datab_exp_not_zero(0);
	wire_w_datab_exp_not_zero_range97w(0) <= datab_exp_not_zero(1);
	wire_w_datab_exp_not_zero_range107w(0) <= datab_exp_not_zero(2);
	wire_w_datab_exp_not_zero_range117w(0) <= datab_exp_not_zero(3);
	wire_w_datab_exp_not_zero_range127w(0) <= datab_exp_not_zero(4);
	wire_w_datab_exp_not_zero_range137w(0) <= datab_exp_not_zero(5);
	wire_w_datab_exp_not_zero_range147w(0) <= datab_exp_not_zero(6);
	wire_w_datab_exp_not_zero_range157w(0) <= datab_exp_not_zero(7);
	wire_w_datab_exp_not_zero_range167w(0) <= datab_exp_not_zero(8);
	wire_w_datab_exp_not_zero_range177w(0) <= datab_exp_not_zero(9);
	wire_w_datab_man_not_zero_range197w(0) <= datab_man_not_zero(0);
	wire_w_datab_man_not_zero_range257w(0) <= datab_man_not_zero(10);
	wire_w_datab_man_not_zero_range263w(0) <= datab_man_not_zero(11);
	wire_w_datab_man_not_zero_range269w(0) <= datab_man_not_zero(12);
	wire_w_datab_man_not_zero_range275w(0) <= datab_man_not_zero(13);
	wire_w_datab_man_not_zero_range281w(0) <= datab_man_not_zero(14);
	wire_w_datab_man_not_zero_range287w(0) <= datab_man_not_zero(15);
	wire_w_datab_man_not_zero_range293w(0) <= datab_man_not_zero(16);
	wire_w_datab_man_not_zero_range299w(0) <= datab_man_not_zero(17);
	wire_w_datab_man_not_zero_range305w(0) <= datab_man_not_zero(18);
	wire_w_datab_man_not_zero_range311w(0) <= datab_man_not_zero(19);
	wire_w_datab_man_not_zero_range203w(0) <= datab_man_not_zero(1);
	wire_w_datab_man_not_zero_range317w(0) <= datab_man_not_zero(20);
	wire_w_datab_man_not_zero_range323w(0) <= datab_man_not_zero(21);
	wire_w_datab_man_not_zero_range329w(0) <= datab_man_not_zero(22);
	wire_w_datab_man_not_zero_range335w(0) <= datab_man_not_zero(23);
	wire_w_datab_man_not_zero_range341w(0) <= datab_man_not_zero(24);
	wire_w_datab_man_not_zero_range352w(0) <= datab_man_not_zero(26);
	wire_w_datab_man_not_zero_range357w(0) <= datab_man_not_zero(27);
	wire_w_datab_man_not_zero_range363w(0) <= datab_man_not_zero(28);
	wire_w_datab_man_not_zero_range369w(0) <= datab_man_not_zero(29);
	wire_w_datab_man_not_zero_range209w(0) <= datab_man_not_zero(2);
	wire_w_datab_man_not_zero_range375w(0) <= datab_man_not_zero(30);
	wire_w_datab_man_not_zero_range381w(0) <= datab_man_not_zero(31);
	wire_w_datab_man_not_zero_range387w(0) <= datab_man_not_zero(32);
	wire_w_datab_man_not_zero_range393w(0) <= datab_man_not_zero(33);
	wire_w_datab_man_not_zero_range399w(0) <= datab_man_not_zero(34);
	wire_w_datab_man_not_zero_range405w(0) <= datab_man_not_zero(35);
	wire_w_datab_man_not_zero_range411w(0) <= datab_man_not_zero(36);
	wire_w_datab_man_not_zero_range417w(0) <= datab_man_not_zero(37);
	wire_w_datab_man_not_zero_range423w(0) <= datab_man_not_zero(38);
	wire_w_datab_man_not_zero_range429w(0) <= datab_man_not_zero(39);
	wire_w_datab_man_not_zero_range215w(0) <= datab_man_not_zero(3);
	wire_w_datab_man_not_zero_range435w(0) <= datab_man_not_zero(40);
	wire_w_datab_man_not_zero_range441w(0) <= datab_man_not_zero(41);
	wire_w_datab_man_not_zero_range447w(0) <= datab_man_not_zero(42);
	wire_w_datab_man_not_zero_range453w(0) <= datab_man_not_zero(43);
	wire_w_datab_man_not_zero_range459w(0) <= datab_man_not_zero(44);
	wire_w_datab_man_not_zero_range465w(0) <= datab_man_not_zero(45);
	wire_w_datab_man_not_zero_range471w(0) <= datab_man_not_zero(46);
	wire_w_datab_man_not_zero_range477w(0) <= datab_man_not_zero(47);
	wire_w_datab_man_not_zero_range483w(0) <= datab_man_not_zero(48);
	wire_w_datab_man_not_zero_range489w(0) <= datab_man_not_zero(49);
	wire_w_datab_man_not_zero_range221w(0) <= datab_man_not_zero(4);
	wire_w_datab_man_not_zero_range495w(0) <= datab_man_not_zero(50);
	wire_w_datab_man_not_zero_range227w(0) <= datab_man_not_zero(5);
	wire_w_datab_man_not_zero_range233w(0) <= datab_man_not_zero(6);
	wire_w_datab_man_not_zero_range239w(0) <= datab_man_not_zero(7);
	wire_w_datab_man_not_zero_range245w(0) <= datab_man_not_zero(8);
	wire_w_datab_man_not_zero_range251w(0) <= datab_man_not_zero(9);
	wire_w_man_result_round_range796w <= man_result_round(50 DOWNTO 0);
	wire_w_man_result_round_range787w(0) <= man_result_round(51);
	wire_w_man_shift_full_range682w <= man_shift_full(53 DOWNTO 1);
	wire_w_result_exp_all_one_range706w(0) <= result_exp_all_one(0);
	wire_w_result_exp_all_one_range709w(0) <= result_exp_all_one(1);
	wire_w_result_exp_all_one_range712w(0) <= result_exp_all_one(2);
	wire_w_result_exp_all_one_range715w(0) <= result_exp_all_one(3);
	wire_w_result_exp_all_one_range718w(0) <= result_exp_all_one(4);
	wire_w_result_exp_all_one_range721w(0) <= result_exp_all_one(5);
	wire_w_result_exp_all_one_range724w(0) <= result_exp_all_one(6);
	wire_w_result_exp_all_one_range727w(0) <= result_exp_all_one(7);
	wire_w_result_exp_all_one_range730w(0) <= result_exp_all_one(8);
	wire_w_result_exp_all_one_range733w(0) <= result_exp_all_one(9);
	wire_w_result_exp_not_zero_range745w(0) <= result_exp_not_zero(0);
	wire_w_result_exp_not_zero_range765w(0) <= result_exp_not_zero(10);
	wire_w_result_exp_not_zero_range767w(0) <= result_exp_not_zero(11);
	wire_w_result_exp_not_zero_range747w(0) <= result_exp_not_zero(1);
	wire_w_result_exp_not_zero_range749w(0) <= result_exp_not_zero(2);
	wire_w_result_exp_not_zero_range751w(0) <= result_exp_not_zero(3);
	wire_w_result_exp_not_zero_range753w(0) <= result_exp_not_zero(4);
	wire_w_result_exp_not_zero_range755w(0) <= result_exp_not_zero(5);
	wire_w_result_exp_not_zero_range757w(0) <= result_exp_not_zero(6);
	wire_w_result_exp_not_zero_range759w(0) <= result_exp_not_zero(7);
	wire_w_result_exp_not_zero_range761w(0) <= result_exp_not_zero(8);
	wire_w_result_exp_not_zero_range763w(0) <= result_exp_not_zero(9);
	wire_w_sticky_bit_range522w(0) <= sticky_bit(0);
	wire_w_sticky_bit_range552w(0) <= sticky_bit(10);
	wire_w_sticky_bit_range555w(0) <= sticky_bit(11);
	wire_w_sticky_bit_range558w(0) <= sticky_bit(12);
	wire_w_sticky_bit_range561w(0) <= sticky_bit(13);
	wire_w_sticky_bit_range564w(0) <= sticky_bit(14);
	wire_w_sticky_bit_range567w(0) <= sticky_bit(15);
	wire_w_sticky_bit_range570w(0) <= sticky_bit(16);
	wire_w_sticky_bit_range573w(0) <= sticky_bit(17);
	wire_w_sticky_bit_range576w(0) <= sticky_bit(18);
	wire_w_sticky_bit_range579w(0) <= sticky_bit(19);
	wire_w_sticky_bit_range525w(0) <= sticky_bit(1);
	wire_w_sticky_bit_range582w(0) <= sticky_bit(20);
	wire_w_sticky_bit_range585w(0) <= sticky_bit(21);
	wire_w_sticky_bit_range588w(0) <= sticky_bit(22);
	wire_w_sticky_bit_range591w(0) <= sticky_bit(23);
	wire_w_sticky_bit_range594w(0) <= sticky_bit(24);
	wire_w_sticky_bit_range597w(0) <= sticky_bit(25);
	wire_w_sticky_bit_range600w(0) <= sticky_bit(26);
	wire_w_sticky_bit_range603w(0) <= sticky_bit(27);
	wire_w_sticky_bit_range606w(0) <= sticky_bit(28);
	wire_w_sticky_bit_range609w(0) <= sticky_bit(29);
	wire_w_sticky_bit_range528w(0) <= sticky_bit(2);
	wire_w_sticky_bit_range612w(0) <= sticky_bit(30);
	wire_w_sticky_bit_range615w(0) <= sticky_bit(31);
	wire_w_sticky_bit_range618w(0) <= sticky_bit(32);
	wire_w_sticky_bit_range621w(0) <= sticky_bit(33);
	wire_w_sticky_bit_range624w(0) <= sticky_bit(34);
	wire_w_sticky_bit_range627w(0) <= sticky_bit(35);
	wire_w_sticky_bit_range630w(0) <= sticky_bit(36);
	wire_w_sticky_bit_range633w(0) <= sticky_bit(37);
	wire_w_sticky_bit_range636w(0) <= sticky_bit(38);
	wire_w_sticky_bit_range639w(0) <= sticky_bit(39);
	wire_w_sticky_bit_range531w(0) <= sticky_bit(3);
	wire_w_sticky_bit_range642w(0) <= sticky_bit(40);
	wire_w_sticky_bit_range645w(0) <= sticky_bit(41);
	wire_w_sticky_bit_range648w(0) <= sticky_bit(42);
	wire_w_sticky_bit_range651w(0) <= sticky_bit(43);
	wire_w_sticky_bit_range654w(0) <= sticky_bit(44);
	wire_w_sticky_bit_range657w(0) <= sticky_bit(45);
	wire_w_sticky_bit_range660w(0) <= sticky_bit(46);
	wire_w_sticky_bit_range663w(0) <= sticky_bit(47);
	wire_w_sticky_bit_range666w(0) <= sticky_bit(48);
	wire_w_sticky_bit_range669w(0) <= sticky_bit(49);
	wire_w_sticky_bit_range534w(0) <= sticky_bit(4);
	wire_w_sticky_bit_range672w(0) <= sticky_bit(50);
	wire_w_sticky_bit_range537w(0) <= sticky_bit(5);
	wire_w_sticky_bit_range540w(0) <= sticky_bit(6);
	wire_w_sticky_bit_range543w(0) <= sticky_bit(7);
	wire_w_sticky_bit_range546w(0) <= sticky_bit(8);
	wire_w_sticky_bit_range549w(0) <= sticky_bit(9);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN dataa_exp_all_one_ff_p1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN dataa_exp_all_one_ff_p1 <= dataa_exp_all_one(10);
			END IF;
		END IF;
	END PROCESS;
	wire_dataa_exp_all_one_ff_p1_w_lg_q512w(0) <= dataa_exp_all_one_ff_p1 AND wire_dataa_man_not_zero_ff_p1_w_lg_w_lg_q506w511w(0);
	wire_dataa_exp_all_one_ff_p1_w_lg_q507w(0) <= dataa_exp_all_one_ff_p1 AND wire_dataa_man_not_zero_ff_p1_w_lg_q506w(0);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN dataa_exp_not_zero_ff_p1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN dataa_exp_not_zero_ff_p1 <= dataa_exp_not_zero(10);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN dataa_man_not_zero_ff_p1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN dataa_man_not_zero_ff_p1 <= dataa_man_not_zero(25);
			END IF;
		END IF;
	END PROCESS;
	wire_dataa_man_not_zero_ff_p1_w_lg_w_lg_q506w511w(0) <= NOT wire_dataa_man_not_zero_ff_p1_w_lg_q506w(0);
	wire_dataa_man_not_zero_ff_p1_w_lg_q506w(0) <= dataa_man_not_zero_ff_p1 OR dataa_man_not_zero_ff_p2;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN dataa_man_not_zero_ff_p2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN dataa_man_not_zero_ff_p2 <= dataa_man_not_zero(51);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN datab_exp_all_one_ff_p1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN datab_exp_all_one_ff_p1 <= datab_exp_all_one(10);
			END IF;
		END IF;
	END PROCESS;
	wire_datab_exp_all_one_ff_p1_w_lg_q510w(0) <= datab_exp_all_one_ff_p1 AND wire_datab_man_not_zero_ff_p1_w_lg_w_lg_q504w509w(0);
	wire_datab_exp_all_one_ff_p1_w_lg_q505w(0) <= datab_exp_all_one_ff_p1 AND wire_datab_man_not_zero_ff_p1_w_lg_q504w(0);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN datab_exp_not_zero_ff_p1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN datab_exp_not_zero_ff_p1 <= datab_exp_not_zero(10);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN datab_man_not_zero_ff_p1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN datab_man_not_zero_ff_p1 <= datab_man_not_zero(25);
			END IF;
		END IF;
	END PROCESS;
	wire_datab_man_not_zero_ff_p1_w_lg_w_lg_q504w509w(0) <= NOT wire_datab_man_not_zero_ff_p1_w_lg_q504w(0);
	wire_datab_man_not_zero_ff_p1_w_lg_q504w(0) <= datab_man_not_zero_ff_p1 OR datab_man_not_zero_ff_p2;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN datab_man_not_zero_ff_p2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN datab_man_not_zero_ff_p2 <= datab_man_not_zero(51);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN delay_exp2_bias <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN delay_exp2_bias <= delay_exp_bias;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN delay_exp_bias <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN delay_exp_bias <= wire_exp_bias_subtr_result;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN delay_man_product_msb <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN delay_man_product_msb <= delay_man_product_msb_p0;
			END IF;
		END IF;
	END PROCESS;
	wire_delay_man_product_msb_w_lg_q696w(0) <= delay_man_product_msb AND wire_man_round_p2_w_q_range694w(0);
	wire_delay_man_product_msb_w_lg_q698w(0) <= delay_man_product_msb XOR wire_man_round_p2_w_q_range694w(0);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN delay_man_product_msb_p0 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN delay_man_product_msb_p0 <= wire_man_product2_mult_w_result_range514w(0);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_add_p1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_add_p1 <= wire_exp_add_adder_result;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_result_ff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_result_ff <= wire_w_lg_w_lg_inf_num777w778w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_dffe_0 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_dffe_0 <= (wire_dataa_exp_all_one_ff_p1_w_lg_q512w(0) OR wire_datab_exp_all_one_ff_p1_w_lg_q510w(0));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_dffe_1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_dffe_1 <= input_is_infinity_dffe_0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_ff1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_ff1 <= input_is_infinity_dffe_1;
			END IF;
		END IF;
	END PROCESS;
	wire_input_is_infinity_ff1_w_lg_q780w(0) <= input_is_infinity_ff1 AND wire_input_not_zero_ff1_w_lg_q779w(0);
	wire_input_is_infinity_ff1_w_lg_q786w(0) <= NOT input_is_infinity_ff1;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_dffe_0 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_dffe_0 <= (wire_dataa_exp_all_one_ff_p1_w_lg_q507w(0) OR wire_datab_exp_all_one_ff_p1_w_lg_q505w(0));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_dffe_1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_dffe_1 <= input_is_nan_dffe_0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_ff1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_ff1 <= input_is_nan_dffe_1;
			END IF;
		END IF;
	END PROCESS;
	wire_input_is_nan_ff1_w_lg_q782w(0) <= NOT input_is_nan_ff1;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_not_zero_dffe_0 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_not_zero_dffe_0 <= (dataa_exp_not_zero_ff_p1 AND datab_exp_not_zero_ff_p1);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_not_zero_dffe_1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_not_zero_dffe_1 <= input_not_zero_dffe_0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_not_zero_ff1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_not_zero_ff1 <= input_not_zero_dffe_1;
			END IF;
		END IF;
	END PROCESS;
	wire_input_not_zero_ff1_w_lg_q779w(0) <= NOT input_not_zero_ff1;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN lsb_dffe <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN lsb_dffe <= lsb_bit;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_result_ff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_result_ff <= ( wire_w_lg_w_lg_w_lg_w790w791w792w793w & wire_w_lg_w_lg_w799w800w801w);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_round_p <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_round_p <= wire_w_man_shift_full_range682w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_round_p2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_round_p2 <= wire_man_round_adder_result;
			END IF;
		END IF;
	END PROCESS;
	loop7 : FOR i IN 0 TO 52 GENERATE 
		wire_man_round_p2_w_lg_w_q_range702w703w(i) <= wire_man_round_p2_w_q_range702w(i) AND wire_man_round_p2_w_lg_w_q_range694w701w(0);
	END GENERATE loop7;
	loop8 : FOR i IN 0 TO 52 GENERATE 
		wire_man_round_p2_w_lg_w_q_range699w700w(i) <= wire_man_round_p2_w_q_range699w(i) AND wire_man_round_p2_w_q_range694w(0);
	END GENERATE loop8;
	wire_man_round_p2_w_lg_w_q_range694w701w(0) <= NOT wire_man_round_p2_w_q_range694w(0);
	wire_man_round_p2_w_q_range702w <= man_round_p2(52 DOWNTO 0);
	wire_man_round_p2_w_q_range699w <= man_round_p2(53 DOWNTO 1);
	wire_man_round_p2_w_q_range694w(0) <= man_round_p2(53);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN overflow_ff <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN overflow_ff <= ((wire_w_lg_exp_is_inf775w(0) AND wire_input_is_nan_ff1_w_lg_q782w(0)) AND (NOT wire_input_is_infinity_ff1_w_lg_q780w(0)));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN round_dffe <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN round_dffe <= round_bit;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_node_ff0 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_node_ff0 <= (dataa(63) XOR datab(63));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_node_ff1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_node_ff1 <= sign_node_ff0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_node_ff2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_node_ff2 <= sign_node_ff1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_node_ff3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_node_ff3 <= sign_node_ff2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_node_ff4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_node_ff4 <= sign_node_ff3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sticky_dffe <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sticky_dffe <= sticky_bit(51);
			END IF;
		END IF;
	END PROCESS;
	wire_exp_add_adder_dataa <= ( "0" & dataa(62 DOWNTO 52));
	wire_exp_add_adder_datab <= ( "0" & datab(62 DOWNTO 52));
	exp_add_adder :  lpm_add_sub
	  GENERIC MAP (
		LPM_PIPELINE => 1,
		LPM_WIDTH => 12
	  )
	  PORT MAP ( 
		aclr => aclr,
		cin => wire_gnd,
		clken => clk_en,
		clock => clock,
		dataa => wire_exp_add_adder_dataa,
		datab => wire_exp_add_adder_datab,
		result => wire_exp_add_adder_result
	  );
	loop9 : FOR i IN 0 TO 10 GENERATE 
		wire_exp_adj_adder_w_lg_w_lg_w_result_range772w773w774w(i) <= wire_exp_adj_adder_w_lg_w_result_range772w773w(i) AND input_not_zero_ff1;
	END GENERATE loop9;
	loop10 : FOR i IN 0 TO 10 GENERATE 
		wire_exp_adj_adder_w_lg_w_result_range772w773w(i) <= wire_exp_adj_adder_w_result_range772w(i) AND wire_w_lg_exp_is_zero771w(0);
	END GENERATE loop10;
	wire_exp_adj_adder_w_lg_w_result_range739w770w(0) <= wire_exp_adj_adder_w_result_range739w(0) OR wire_w_lg_w_result_exp_not_zero_range767w769w(0);
	wire_exp_adj_adder_w_result_range772w <= wire_exp_adj_adder_result(10 DOWNTO 0);
	wire_exp_adj_adder_w_result_range735w(0) <= wire_exp_adj_adder_result(10);
	wire_exp_adj_adder_w_result_range738w(0) <= wire_exp_adj_adder_result(11);
	wire_exp_adj_adder_w_result_range739w(0) <= wire_exp_adj_adder_result(12);
	wire_exp_adj_adder_w_result_range708w(0) <= wire_exp_adj_adder_result(1);
	wire_exp_adj_adder_w_result_range711w(0) <= wire_exp_adj_adder_result(2);
	wire_exp_adj_adder_w_result_range714w(0) <= wire_exp_adj_adder_result(3);
	wire_exp_adj_adder_w_result_range717w(0) <= wire_exp_adj_adder_result(4);
	wire_exp_adj_adder_w_result_range720w(0) <= wire_exp_adj_adder_result(5);
	wire_exp_adj_adder_w_result_range723w(0) <= wire_exp_adj_adder_result(6);
	wire_exp_adj_adder_w_result_range726w(0) <= wire_exp_adj_adder_result(7);
	wire_exp_adj_adder_w_result_range729w(0) <= wire_exp_adj_adder_result(8);
	wire_exp_adj_adder_w_result_range732w(0) <= wire_exp_adj_adder_result(9);
	exp_adj_adder :  lpm_add_sub
	  GENERIC MAP (
		LPM_WIDTH => 13
	  )
	  PORT MAP ( 
		cin => wire_gnd,
		dataa => delay_exp2_bias,
		datab => expmod,
		result => wire_exp_adj_adder_result
	  );
	wire_exp_bias_subtr_dataa <= ( "0" & exp_add_p1(11 DOWNTO 0));
	wire_exp_bias_subtr_datab <= ( bias(12 DOWNTO 0));
	exp_bias_subtr :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_PIPELINE => 0,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 13
	  )
	  PORT MAP ( 
		dataa => wire_exp_bias_subtr_dataa,
		datab => wire_exp_bias_subtr_datab,
		result => wire_exp_bias_subtr_result
	  );
	wire_man_round_adder_dataa <= ( "0" & man_round_p);
	wire_man_round_adder_datab <= ( "00000000000000000000000000000000000000000000000000000" & round_carry);
	man_round_adder :  lpm_add_sub
	  GENERIC MAP (
		LPM_PIPELINE => 0,
		LPM_WIDTH => 54
	  )
	  PORT MAP ( 
		dataa => wire_man_round_adder_dataa,
		datab => wire_man_round_adder_datab,
		result => wire_man_round_adder_result
	  );
	loop11 : FOR i IN 0 TO 53 GENERATE 
		wire_man_product2_mult_w_lg_w_result_range518w519w(i) <= wire_man_product2_mult_w_result_range518w(i) AND wire_man_product2_mult_w_lg_w_result_range514w517w(0);
	END GENERATE loop11;
	wire_man_product2_mult_w_lg_w_result_range514w676w(0) <= wire_man_product2_mult_w_result_range514w(0) AND wire_man_product2_mult_w_result_range674w(0);
	loop12 : FOR i IN 0 TO 53 GENERATE 
		wire_man_product2_mult_w_lg_w_result_range515w516w(i) <= wire_man_product2_mult_w_result_range515w(i) AND wire_man_product2_mult_w_result_range514w(0);
	END GENERATE loop12;
	wire_man_product2_mult_w_lg_w_result_range514w517w(0) <= NOT wire_man_product2_mult_w_result_range514w(0);
	wire_man_product2_mult_dataa <= ( "1" & dataa(51 DOWNTO 0));
	wire_man_product2_mult_datab <= ( "1" & datab(51 DOWNTO 0));
	wire_man_product2_mult_w_result_range518w <= wire_man_product2_mult_result(104 DOWNTO 51);
	wire_man_product2_mult_w_result_range514w(0) <= wire_man_product2_mult_result(105);
	wire_man_product2_mult_w_result_range515w <= wire_man_product2_mult_result(105 DOWNTO 52);
	wire_man_product2_mult_w_result_range551w(0) <= wire_man_product2_mult_result(10);
	wire_man_product2_mult_w_result_range554w(0) <= wire_man_product2_mult_result(11);
	wire_man_product2_mult_w_result_range557w(0) <= wire_man_product2_mult_result(12);
	wire_man_product2_mult_w_result_range560w(0) <= wire_man_product2_mult_result(13);
	wire_man_product2_mult_w_result_range563w(0) <= wire_man_product2_mult_result(14);
	wire_man_product2_mult_w_result_range566w(0) <= wire_man_product2_mult_result(15);
	wire_man_product2_mult_w_result_range569w(0) <= wire_man_product2_mult_result(16);
	wire_man_product2_mult_w_result_range572w(0) <= wire_man_product2_mult_result(17);
	wire_man_product2_mult_w_result_range575w(0) <= wire_man_product2_mult_result(18);
	wire_man_product2_mult_w_result_range578w(0) <= wire_man_product2_mult_result(19);
	wire_man_product2_mult_w_result_range524w(0) <= wire_man_product2_mult_result(1);
	wire_man_product2_mult_w_result_range581w(0) <= wire_man_product2_mult_result(20);
	wire_man_product2_mult_w_result_range584w(0) <= wire_man_product2_mult_result(21);
	wire_man_product2_mult_w_result_range587w(0) <= wire_man_product2_mult_result(22);
	wire_man_product2_mult_w_result_range590w(0) <= wire_man_product2_mult_result(23);
	wire_man_product2_mult_w_result_range593w(0) <= wire_man_product2_mult_result(24);
	wire_man_product2_mult_w_result_range596w(0) <= wire_man_product2_mult_result(25);
	wire_man_product2_mult_w_result_range599w(0) <= wire_man_product2_mult_result(26);
	wire_man_product2_mult_w_result_range602w(0) <= wire_man_product2_mult_result(27);
	wire_man_product2_mult_w_result_range605w(0) <= wire_man_product2_mult_result(28);
	wire_man_product2_mult_w_result_range608w(0) <= wire_man_product2_mult_result(29);
	wire_man_product2_mult_w_result_range527w(0) <= wire_man_product2_mult_result(2);
	wire_man_product2_mult_w_result_range611w(0) <= wire_man_product2_mult_result(30);
	wire_man_product2_mult_w_result_range614w(0) <= wire_man_product2_mult_result(31);
	wire_man_product2_mult_w_result_range617w(0) <= wire_man_product2_mult_result(32);
	wire_man_product2_mult_w_result_range620w(0) <= wire_man_product2_mult_result(33);
	wire_man_product2_mult_w_result_range623w(0) <= wire_man_product2_mult_result(34);
	wire_man_product2_mult_w_result_range626w(0) <= wire_man_product2_mult_result(35);
	wire_man_product2_mult_w_result_range629w(0) <= wire_man_product2_mult_result(36);
	wire_man_product2_mult_w_result_range632w(0) <= wire_man_product2_mult_result(37);
	wire_man_product2_mult_w_result_range635w(0) <= wire_man_product2_mult_result(38);
	wire_man_product2_mult_w_result_range638w(0) <= wire_man_product2_mult_result(39);
	wire_man_product2_mult_w_result_range530w(0) <= wire_man_product2_mult_result(3);
	wire_man_product2_mult_w_result_range641w(0) <= wire_man_product2_mult_result(40);
	wire_man_product2_mult_w_result_range644w(0) <= wire_man_product2_mult_result(41);
	wire_man_product2_mult_w_result_range647w(0) <= wire_man_product2_mult_result(42);
	wire_man_product2_mult_w_result_range650w(0) <= wire_man_product2_mult_result(43);
	wire_man_product2_mult_w_result_range653w(0) <= wire_man_product2_mult_result(44);
	wire_man_product2_mult_w_result_range656w(0) <= wire_man_product2_mult_result(45);
	wire_man_product2_mult_w_result_range659w(0) <= wire_man_product2_mult_result(46);
	wire_man_product2_mult_w_result_range662w(0) <= wire_man_product2_mult_result(47);
	wire_man_product2_mult_w_result_range665w(0) <= wire_man_product2_mult_result(48);
	wire_man_product2_mult_w_result_range668w(0) <= wire_man_product2_mult_result(49);
	wire_man_product2_mult_w_result_range533w(0) <= wire_man_product2_mult_result(4);
	wire_man_product2_mult_w_result_range671w(0) <= wire_man_product2_mult_result(50);
	wire_man_product2_mult_w_result_range674w(0) <= wire_man_product2_mult_result(51);
	wire_man_product2_mult_w_result_range536w(0) <= wire_man_product2_mult_result(5);
	wire_man_product2_mult_w_result_range539w(0) <= wire_man_product2_mult_result(6);
	wire_man_product2_mult_w_result_range542w(0) <= wire_man_product2_mult_result(7);
	wire_man_product2_mult_w_result_range545w(0) <= wire_man_product2_mult_result(8);
	wire_man_product2_mult_w_result_range548w(0) <= wire_man_product2_mult_result(9);
	man_product2_mult :  lpm_mult
	  GENERIC MAP (
		LPM_PIPELINE => 2,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTHA => 53,
		LPM_WIDTHB => 53,
		LPM_WIDTHP => 106,
		LPM_WIDTHS => 1,
		lpm_hint => "DEDICATED_MULTIPLIER_CIRCUITRY=YES"
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => wire_man_product2_mult_dataa,
		datab => wire_man_product2_mult_datab,
		result => wire_man_product2_mult_result
	  );

 END RTL; --mult_altfp_mult_nto
--VALID FILE


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY mult IS
	PORT
	(
		clock		: IN STD_LOGIC ;
		dataa		: IN STD_LOGIC_VECTOR (63 DOWNTO 0);
		datab		: IN STD_LOGIC_VECTOR (63 DOWNTO 0);
		overflow		: OUT STD_LOGIC ;
		result		: OUT STD_LOGIC_VECTOR (63 DOWNTO 0)
	);
END mult;


ARCHITECTURE RTL OF mult IS

	SIGNAL sub_wire0	: STD_LOGIC ;
	SIGNAL sub_wire1	: STD_LOGIC_VECTOR (63 DOWNTO 0);



	COMPONENT mult_altfp_mult_nto
	PORT (
			clock	: IN STD_LOGIC ;
			datab	: IN STD_LOGIC_VECTOR (63 DOWNTO 0);
			overflow	: OUT STD_LOGIC ;
			dataa	: IN STD_LOGIC_VECTOR (63 DOWNTO 0);
			result	: OUT STD_LOGIC_VECTOR (63 DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	overflow    <= sub_wire0;
	result    <= sub_wire1(63 DOWNTO 0);

	mult_altfp_mult_nto_component : mult_altfp_mult_nto
	PORT MAP (
		clock => clock,
		datab => datab,
		dataa => dataa,
		overflow => sub_wire0,
		result => sub_wire1
	);



END RTL;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: PRIVATE: FPM_FORMAT STRING "Double"
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone IV GX"
-- Retrieval info: CONSTANT: DEDICATED_MULTIPLIER_CIRCUITRY STRING "YES"
-- Retrieval info: CONSTANT: DENORMAL_SUPPORT STRING "NO"
-- Retrieval info: CONSTANT: EXCEPTION_HANDLING STRING "NO"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "UNUSED"
-- Retrieval info: CONSTANT: LPM_HINT STRING "UNUSED"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "altfp_mult"
-- Retrieval info: CONSTANT: PIPELINE NUMERIC "5"
-- Retrieval info: CONSTANT: REDUCED_FUNCTIONALITY STRING "NO"
-- Retrieval info: CONSTANT: ROUNDING STRING "TO_NEAREST"
-- Retrieval info: CONSTANT: WIDTH_EXP NUMERIC "11"
-- Retrieval info: CONSTANT: WIDTH_MAN NUMERIC "52"
-- Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL "clock"
-- Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
-- Retrieval info: USED_PORT: dataa 0 0 64 0 INPUT NODEFVAL "dataa[63..0]"
-- Retrieval info: CONNECT: @dataa 0 0 64 0 dataa 0 0 64 0
-- Retrieval info: USED_PORT: datab 0 0 64 0 INPUT NODEFVAL "datab[63..0]"
-- Retrieval info: CONNECT: @datab 0 0 64 0 datab 0 0 64 0
-- Retrieval info: USED_PORT: overflow 0 0 0 0 OUTPUT NODEFVAL "overflow"
-- Retrieval info: CONNECT: overflow 0 0 0 0 @overflow 0 0 0 0
-- Retrieval info: USED_PORT: result 0 0 64 0 OUTPUT NODEFVAL "result[63..0]"
-- Retrieval info: CONNECT: result 0 0 64 0 @result 0 0 64 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL mult.vhd TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL mult.qip TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL mult.bsf TRUE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL mult_inst.vhd TRUE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL mult.inc TRUE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL mult.cmp TRUE TRUE
-- Retrieval info: LIB_FILE: lpm
